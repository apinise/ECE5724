module c5315_tb (
);

reg [1:178] n;
wire [122:0] o, onet;

c5315 GUT (
  // Inputs
  .N1(n[1]),
  .N4(n[2]),
  .N11(n[3]),
  .N14(n[4]),
  .N17(n[5]),
  .N20(n[6]),
  .N23(n[7]),
  .N24(n[8]),
  .N25(n[9]),
  .N26(n[10]),
  .N27(n[11]),
  .N31(n[12]),
  .N34(n[13]),
  .N37(n[14]),
  .N40(n[15]),
  .N43(n[16]),
  .N46(n[17]),
  .N49(n[18]),
  .N52(n[19]),
  .N53(n[20]),
  .N54(n[21]),
  .N61(n[22]),
  .N64(n[23]),
  .N67(n[24]),
  .N70(n[25]),
  .N73(n[26]),
  .N76(n[27]),
  .N79(n[28]),
  .N80(n[29]),
  .N81(n[30]),
  .N82(n[31]),
  .N83(n[32]),
  .N86(n[33]),
  .N87(n[34]),
  .N88(n[35]),
  .N91(n[36]),
  .N94(n[37]),
  .N97(n[38]),
  .N100(n[39]),
  .N103(n[40]),
  .N106(n[41]),
  .N109(n[42]),
  .N112(n[43]),
  .N113(n[44]),
  .N114(n[45]),
  .N115(n[46]),
  .N116(n[47]),
  .N117(n[48]),
  .N118(n[49]),
  .N119(n[50]),
  .N120(n[51]),
  .N121(n[52]),
  .N122(n[53]),
  .N123(n[54]),
  .N126(n[55]),
  .N127(n[56]),
  .N128(n[57]),
  .N129(n[58]),
  .N130(n[59]),
  .N131(n[60]),
  .N132(n[61]),
  .N135(n[62]),
  .N136(n[63]),
  .N137(n[64]),
  .N140(n[65]),
  .N141(n[66]),
  .N145(n[67]),
  .N146(n[68]),
  .N149(n[69]),
  .N152(n[70]),
  .N155(n[71]),
  .N158(n[72]),
  .N161(n[73]),
  .N164(n[74]),
  .N167(n[75]),
  .N170(n[76]),
  .N173(n[77]),
  .N176(n[78]),
  .N179(n[79]),
  .N182(n[80]),
  .N185(n[81]),
  .N188(n[82]),
  .N191(n[83]),
  .N194(n[84]),
  .N197(n[85]),
  .N200(n[86]),
  .N203(n[87]),
  .N206(n[88]),
  .N209(n[89]),
  .N210(n[90]),
  .N217(n[91]),
  .N218(),
  .N225(),
  .N226(),
  .N233(),
  .N234(),
  .N241(),
  .N242(),
  .N245(),
  .N248(),
  .N251(),
  .N254(),
  .N257(),
  .N264(),
  .N265(),
  .N272(),
  .N273(),
  .N280(),
  .N281(),
  .N288(),
  .N289(),
  .N292(),
  .N293(),
  .N299(),
  .N302(),
  .N307(),
  .N308(),
  .N315(),
  .N316(),
  .N323(),
  .N324(),
  .N331(),
  .N332(),
  .N335(),
  .N338(),
  .N341(),
  .N348(),
  .N351(),
  .N358(),
  .N361(),
  .N366(),
  .N369(),
  .N372(),
  .N373(),
  .N374(),
  .N386(),
  .N389(),
  .N400(),
  .N411(),
  .N422(),
  .N435(),
  .N446(),
  .N457(),
  .N468(),
  .N479(),
  .N490(),
  .N503(),
  .N514(),
  .N523(),
  .N534(),
  .N545(),
  .N549(),
  .N552(),
  .N556(),
  .N559(),
  .N562(),
  .N566(),
  .N571(),
  .N574(),
  .N577(),
  .N580(),
  .N583(),
  .N588(),
  .N591(),
  .N592(),
  .N595(),
  .N596(),
  .N597(),
  .N598(),
  .N599(),
  .N603(),
  .N607(),
  .N610(),
  .N613(),
  .N616(),
  .N619(),
  .N625(),
  .N631(),
  // Outputs
  .N709(),
  .N816(),
  .N1066(),
  .N1137(),
  .N1138(),
  .N1139(),
  .N1140(),
  .N1141(),
  .N1142(),
  .N1143(),
  .N1144(),
  .N1145(),
  .N1147(),
  .N1152(),
  .N1153(),
  .N1154(),
  .N1155(),
  .N1972(),
  .N2054(),
  .N2060(),
  .N2061(),
  .N2139(),
  .N2142(),
  .N2309(),
  .N2387(),
  .N2527(),
  .N2584(),
  .N2590(),
  .N2623(),
  .N3357(),
  .N3358(),
  .N3359(),
  .N3360(),
  .N3604(),
  .N3613(),
  .N4272(),
  .N4275(),
  .N4278(),
  .N4279(),
  .N4737(),
  .N4738(),
  .N4739(),
  .N4740(),
  .N5240(),
  .N5388(),
  .N6641(),
  .N6643(),
  .N6646(),
  .N6648(),
  .N6716(),
  .N6877(),
  .N6924(),
  .N6925(),
  .N6926(),
  .N6927(),
  .N7015(),
  .N7363(),
  .N7365(),
  .N7432(),
  .N7449(),
  .N7465(),
  .N7466(),
  .N7467(),
  .N7469(),
  .N7470(),
  .N7471(),
  .N7472(),
  .N7473(),
  .N7474(),
  .N7476(),
  .N7503(),
  .N7504(),
  .N7506(),
  .N7511(),
  .N7515(),
  .N7516(),
  .N7517(),
  .N7518(),
  .N7519(),
  .N7520(),
  .N7521(),
  .N7522(),
  .N7600(),
  .N7601(),
  .N7602(),
  .N7603(),
  .N7604(),
  .N7605(),
  .N7606(),
  .N7607(),
  .N7626(),
  .N7698(),
  .N7699(),
  .N7700(),
  .N7701(),
  .N7702(),
  .N7703(),
  .N7704(),
  .N7705(),
  .N7706(),
  .N7707(),
  .N7735(),
  .N7736(),
  .N7737(),
  .N7738(),
  .N7739(),
  .N7740(),
  .N7741(),
  .N7742(),
  .N7754(),
  .N7755(),
  .N7756(),
  .N7757(),
  .N7758(),
  .N7759(),
  .N7760(),
  .N7761(),
  .N8075(),
  .N8076(),
  .N8123(),
  .N8124(),
  .N8127(),
  .N8128()
);

endmodule