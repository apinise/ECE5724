`timescale 1ns / 1ps

module c5315_tb (
);

parameter numOfFault = 5104;
parameter inputWidth = 178;
parameter outputWidth = 123;
parameter initialExpFCount = 2; 
parameter utLimit = 20; 
parameter desiredCoverage = 90; 

reg [1:inputWidth] n;
wire [outputWidth-1:0] o, onet;

reg detected = 0;
integer i;
integer faultFile, testFile, status; 
integer uTests, detectedFaultsCT, expFCountCT, faultIndex; 
integer tmp, newDiscovered, coverage, detectedFaultsAT; 
integer keepedCT, totalCT;
real numOfFaults = 5104;
real numOfDetecteds = 0;
real coverage = 0;
reg[1:inputWidth] testVector;
reg[60*8:1] wireName;
reg stuckAtVal;
reg [1:numOfFaults] detectedListCT, detectedListAT;


c5315_net GUT (
  // Inputs
  .N1(n[1]),
  .N4(n[2]),
  .N11(n[3]),
  .N14(n[4]),
  .N17(n[5]),
  .N20(n[6]),
  .N23(n[7]),
  .N24(n[8]),
  .N25(n[9]),
  .N26(n[10]),
  .N27(n[11]),
  .N31(n[12]),
  .N34(n[13]),
  .N37(n[14]),
  .N40(n[15]),
  .N43(n[16]),
  .N46(n[17]),
  .N49(n[18]),
  .N52(n[19]),
  .N53(n[20]),
  .N54(n[21]),
  .N61(n[22]),
  .N64(n[23]),
  .N67(n[24]),
  .N70(n[25]),
  .N73(n[26]),
  .N76(n[27]),
  .N79(n[28]),
  .N80(n[29]),
  .N81(n[30]),
  .N82(n[31]),
  .N83(n[32]),
  .N86(n[33]),
  .N87(n[34]),
  .N88(n[35]),
  .N91(n[36]),
  .N94(n[37]),
  .N97(n[38]),
  .N100(n[39]),
  .N103(n[40]),
  .N106(n[41]),
  .N109(n[42]),
  .N112(n[43]),
  .N113(n[44]),
  .N114(n[45]),
  .N115(n[46]),
  .N116(n[47]),
  .N117(n[48]),
  .N118(n[49]),
  .N119(n[50]),
  .N120(n[51]),
  .N121(n[52]),
  .N122(n[53]),
  .N123(n[54]),
  .N126(n[55]),
  .N127(n[56]),
  .N128(n[57]),
  .N129(n[58]),
  .N130(n[59]),
  .N131(n[60]),
  .N132(n[61]),
  .N135(n[62]),
  .N136(n[63]),
  .N137(n[64]),
  .N140(n[65]),
  .N141(n[66]),
  .N145(n[67]),
  .N146(n[68]),
  .N149(n[69]),
  .N152(n[70]),
  .N155(n[71]),
  .N158(n[72]),
  .N161(n[73]),
  .N164(n[74]),
  .N167(n[75]),
  .N170(n[76]),
  .N173(n[77]),
  .N176(n[78]),
  .N179(n[79]),
  .N182(n[80]),
  .N185(n[81]),
  .N188(n[82]),
  .N191(n[83]),
  .N194(n[84]),
  .N197(n[85]),
  .N200(n[86]),
  .N203(n[87]),
  .N206(n[88]),
  .N209(n[89]),
  .N210(n[90]),
  .N217(n[91]),
  .N218(n[92]),
  .N225(n[93]),
  .N226(n[94]),
  .N233(n[95]),
  .N234(n[96]),
  .N241(n[97]),
  .N242(n[98]),
  .N245(n[99]),
  .N248(n[100]),
  .N251(n[101]),
  .N254(n[102]),
  .N257(n[103]),
  .N264(n[104]),
  .N265(n[105]),
  .N272(n[106]),
  .N273(n[107]),
  .N280(n[108]),
  .N281(n[109]),
  .N288(n[110]),
  .N289(n[111]),
  .N292(n[112]),
  .N293(n[113]),
  .N299(n[114]),
  .N302(n[115]),
  .N307(n[116]),
  .N308(n[117]),
  .N315(n[118]),
  .N316(n[119]),
  .N323(n[120]),
  .N324(n[121]),
  .N331(n[122]),
  .N332(n[123]),
  .N335(n[124]),
  .N338(n[125]),
  .N341(n[126]),
  .N348(n[127]),
  .N351(n[128]),
  .N358(n[129]),
  .N361(n[130]),
  .N366(n[131]),
  .N369(n[132]),
  .N372(n[133]),
  .N373(n[134]),
  .N374(n[135]),
  .N386(n[136]),
  .N389(n[137]),
  .N400(n[138]),
  .N411(n[139]),
  .N422(n[140]),
  .N435(n[141]),
  .N446(n[142]),
  .N457(n[143]),
  .N468(n[144]),
  .N479(n[145]),
  .N490(n[146]),
  .N503(n[147]),
  .N514(n[148]),
  .N523(n[149]),
  .N534(n[150]),
  .N545(n[151]),
  .N549(n[152]),
  .N552(n[153]),
  .N556(n[154]),
  .N559(n[155]),
  .N562(n[156]),
  .N566(n[157]),
  .N571(n[158]),
  .N574(n[159]),
  .N577(n[160]),
  .N580(n[161]),
  .N583(n[162]),
  .N588(n[163]),
  .N591(n[164]),
  .N592(n[165]),
  .N595(n[166]),
  .N596(n[167]),
  .N597(n[168]),
  .N598(n[169]),
  .N599(n[170]),
  .N603(n[171]),
  .N607(n[172]),
  .N610(n[173]),
  .N613(n[174]),
  .N616(n[175]),
  .N619(n[176]),
  .N625(n[177]),
  .N631(n[178]),
  // Outputs
  .N709(o[0]),
  .N816(o[1]),
  .N1066(o[2]),
  .N1137(o[3]),
  .N1138(o[4]),
  .N1139(o[5]),
  .N1140(o[6]),
  .N1141(o[7]),
  .N1142(o[8]),
  .N1143(o[9]),
  .N1144(o[10]),
  .N1145(o[11]),
  .N1147(o[12]),
  .N1152(o[13]),
  .N1153(o[14]),
  .N1154(o[15]),
  .N1155(o[16]),
  .N1972(o[17]),
  .N2054(o[18]),
  .N2060(o[19]),
  .N2061(o[20]),
  .N2139(o[21]),
  .N2142(o[22]),
  .N2309(o[23]),
  .N2387(o[24]),
  .N2527(o[25]),
  .N2584(o[26]),
  .N2590(o[27]),
  .N2623(o[28]),
  .N3357(o[29]),
  .N3358(o[30]),
  .N3359(o[31]),
  .N3360(o[32]),
  .N3604(o[33]),
  .N3613(o[34]),
  .N4272(o[35]),
  .N4275(o[36]),
  .N4278(o[37]),
  .N4279(o[38]),
  .N4737(o[39]),
  .N4738(o[40]),
  .N4739(o[41]),
  .N4740(o[42]),
  .N5240(o[43]),
  .N5388(o[44]),
  .N6641(o[45]),
  .N6643(o[46]),
  .N6646(o[47]),
  .N6648(o[48]),
  .N6716(o[49]),
  .N6877(o[50]),
  .N6924(o[51]),
  .N6925(o[52]),
  .N6926(o[53]),
  .N6927(o[54]),
  .N7015(o[55]),
  .N7363(o[56]),
  .N7365(o[57]),
  .N7432(o[58]),
  .N7449(o[59]),
  .N7465(o[60]),
  .N7466(o[61]),
  .N7467(o[62]),
  .N7469(o[63]),
  .N7470(o[64]),
  .N7471(o[65]),
  .N7472(o[66]),
  .N7473(o[67]),
  .N7474(o[68]),
  .N7476(o[69]),
  .N7503(o[70]),
  .N7504(o[71]),
  .N7506(o[72]),
  .N7511(o[73]),
  .N7515(o[74]),
  .N7516(o[75]),
  .N7517(o[76]),
  .N7518(o[77]),
  .N7519(o[78]),
  .N7520(o[79]),
  .N7521(o[80]),
  .N7522(o[81]),
  .N7600(o[82]),
  .N7601(o[83]),
  .N7602(o[84]),
  .N7603(o[85]),
  .N7604(o[86]),
  .N7605(o[87]),
  .N7606(o[88]),
  .N7607(o[89]),
  .N7626(o[90]),
  .N7698(o[91]),
  .N7699(o[92]),
  .N7700(o[93]),
  .N7701(o[94]),
  .N7702(o[95]),
  .N7703(o[96]),
  .N7704(o[97]),
  .N7705(o[98]),
  .N7706(o[99]),
  .N7707(o[100]),
  .N7735(o[101]),
  .N7736(o[102]),
  .N7737(o[103]),
  .N7738(o[104]),
  .N7739(o[105]),
  .N7740(o[106]),
  .N7741(o[107]),
  .N7742(o[108]),
  .N7754(o[109]),
  .N7755(o[110]),
  .N7756(o[111]),
  .N7757(o[112]),
  .N7758(o[113]),
  .N7759(o[114]),
  .N7760(o[115]),
  .N7761(o[116]),
  .N8075(o[117]),
  .N8076(o[118]),
  .N8123(o[119]),
  .N8124(o[120]),
  .N8127(o[121]),
  .N8128(o[122])
);

c5315_net FUT (
  // Inputs
  .N1(n[1]),
  .N4(n[2]),
  .N11(n[3]),
  .N14(n[4]),
  .N17(n[5]),
  .N20(n[6]),
  .N23(n[7]),
  .N24(n[8]),
  .N25(n[9]),
  .N26(n[10]),
  .N27(n[11]),
  .N31(n[12]),
  .N34(n[13]),
  .N37(n[14]),
  .N40(n[15]),
  .N43(n[16]),
  .N46(n[17]),
  .N49(n[18]),
  .N52(n[19]),
  .N53(n[20]),
  .N54(n[21]),
  .N61(n[22]),
  .N64(n[23]),
  .N67(n[24]),
  .N70(n[25]),
  .N73(n[26]),
  .N76(n[27]),
  .N79(n[28]),
  .N80(n[29]),
  .N81(n[30]),
  .N82(n[31]),
  .N83(n[32]),
  .N86(n[33]),
  .N87(n[34]),
  .N88(n[35]),
  .N91(n[36]),
  .N94(n[37]),
  .N97(n[38]),
  .N100(n[39]),
  .N103(n[40]),
  .N106(n[41]),
  .N109(n[42]),
  .N112(n[43]),
  .N113(n[44]),
  .N114(n[45]),
  .N115(n[46]),
  .N116(n[47]),
  .N117(n[48]),
  .N118(n[49]),
  .N119(n[50]),
  .N120(n[51]),
  .N121(n[52]),
  .N122(n[53]),
  .N123(n[54]),
  .N126(n[55]),
  .N127(n[56]),
  .N128(n[57]),
  .N129(n[58]),
  .N130(n[59]),
  .N131(n[60]),
  .N132(n[61]),
  .N135(n[62]),
  .N136(n[63]),
  .N137(n[64]),
  .N140(n[65]),
  .N141(n[66]),
  .N145(n[67]),
  .N146(n[68]),
  .N149(n[69]),
  .N152(n[70]),
  .N155(n[71]),
  .N158(n[72]),
  .N161(n[73]),
  .N164(n[74]),
  .N167(n[75]),
  .N170(n[76]),
  .N173(n[77]),
  .N176(n[78]),
  .N179(n[79]),
  .N182(n[80]),
  .N185(n[81]),
  .N188(n[82]),
  .N191(n[83]),
  .N194(n[84]),
  .N197(n[85]),
  .N200(n[86]),
  .N203(n[87]),
  .N206(n[88]),
  .N209(n[89]),
  .N210(n[90]),
  .N217(n[91]),
  .N218(n[92]),
  .N225(n[93]),
  .N226(n[94]),
  .N233(n[95]),
  .N234(n[96]),
  .N241(n[97]),
  .N242(n[98]),
  .N245(n[99]),
  .N248(n[100]),
  .N251(n[101]),
  .N254(n[102]),
  .N257(n[103]),
  .N264(n[104]),
  .N265(n[105]),
  .N272(n[106]),
  .N273(n[107]),
  .N280(n[108]),
  .N281(n[109]),
  .N288(n[110]),
  .N289(n[111]),
  .N292(n[112]),
  .N293(n[113]),
  .N299(n[114]),
  .N302(n[115]),
  .N307(n[116]),
  .N308(n[117]),
  .N315(n[118]),
  .N316(n[119]),
  .N323(n[120]),
  .N324(n[121]),
  .N331(n[122]),
  .N332(n[123]),
  .N335(n[124]),
  .N338(n[125]),
  .N341(n[126]),
  .N348(n[127]),
  .N351(n[128]),
  .N358(n[129]),
  .N361(n[130]),
  .N366(n[131]),
  .N369(n[132]),
  .N372(n[133]),
  .N373(n[134]),
  .N374(n[135]),
  .N386(n[136]),
  .N389(n[137]),
  .N400(n[138]),
  .N411(n[139]),
  .N422(n[140]),
  .N435(n[141]),
  .N446(n[142]),
  .N457(n[143]),
  .N468(n[144]),
  .N479(n[145]),
  .N490(n[146]),
  .N503(n[147]),
  .N514(n[148]),
  .N523(n[149]),
  .N534(n[150]),
  .N545(n[151]),
  .N549(n[152]),
  .N552(n[153]),
  .N556(n[154]),
  .N559(n[155]),
  .N562(n[156]),
  .N566(n[157]),
  .N571(n[158]),
  .N574(n[159]),
  .N577(n[160]),
  .N580(n[161]),
  .N583(n[162]),
  .N588(n[163]),
  .N591(n[164]),
  .N592(n[165]),
  .N595(n[166]),
  .N596(n[167]),
  .N597(n[168]),
  .N598(n[169]),
  .N599(n[170]),
  .N603(n[171]),
  .N607(n[172]),
  .N610(n[173]),
  .N613(n[174]),
  .N616(n[175]),
  .N619(n[176]),
  .N625(n[177]),
  .N631(n[178]),
  // Outputs
  .N709(onet[0]),
  .N816(onet[1]),
  .N1066(onet[2]),
  .N1137(onet[3]),
  .N1138(onet[4]),
  .N1139(onet[5]),
  .N1140(onet[6]),
  .N1141(onet[7]),
  .N1142(onet[8]),
  .N1143(onet[9]),
  .N1144(onet[10]),
  .N1145(onet[11]),
  .N1147(onet[12]),
  .N1152(onet[13]),
  .N1153(onet[14]),
  .N1154(onet[15]),
  .N1155(onet[16]),
  .N1972(onet[17]),
  .N2054(onet[18]),
  .N2060(onet[19]),
  .N2061(onet[20]),
  .N2139(onet[21]),
  .N2142(onet[22]),
  .N2309(onet[23]),
  .N2387(onet[24]),
  .N2527(onet[25]),
  .N2584(onet[26]),
  .N2590(onet[27]),
  .N2623(onet[28]),
  .N3357(onet[29]),
  .N3358(onet[30]),
  .N3359(onet[31]),
  .N3360(onet[32]),
  .N3604(onet[33]),
  .N3613(onet[34]),
  .N4272(onet[35]),
  .N4275(onet[36]),
  .N4278(onet[37]),
  .N4279(onet[38]),
  .N4737(onet[39]),
  .N4738(onet[40]),
  .N4739(onet[41]),
  .N4740(onet[42]),
  .N5240(onet[43]),
  .N5388(onet[44]),
  .N6641(onet[45]),
  .N6643(onet[46]),
  .N6646(onet[47]),
  .N6648(onet[48]),
  .N6716(onet[49]),
  .N6877(onet[50]),
  .N6924(onet[51]),
  .N6925(onet[52]),
  .N6926(onet[53]),
  .N6927(onet[54]),
  .N7015(onet[55]),
  .N7363(onet[56]),
  .N7365(onet[57]),
  .N7432(onet[58]),
  .N7449(onet[59]),
  .N7465(onet[60]),
  .N7466(onet[61]),
  .N7467(onet[62]),
  .N7469(onet[63]),
  .N7470(onet[64]),
  .N7471(onet[65]),
  .N7472(onet[66]),
  .N7473(onet[67]),
  .N7474(onet[68]),
  .N7476(onet[69]),
  .N7503(onet[70]),
  .N7504(onet[71]),
  .N7506(onet[72]),
  .N7511(onet[73]),
  .N7515(onet[74]),
  .N7516(onet[75]),
  .N7517(onet[76]),
  .N7518(onet[77]),
  .N7519(onet[78]),
  .N7520(onet[79]),
  .N7521(onet[80]),
  .N7522(onet[81]),
  .N7600(onet[82]),
  .N7601(onet[83]),
  .N7602(onet[84]),
  .N7603(onet[85]),
  .N7604(onet[86]),
  .N7605(onet[87]),
  .N7606(onet[88]),
  .N7607(onet[89]),
  .N7626(onet[90]),
  .N7698(onet[91]),
  .N7699(onet[92]),
  .N7700(onet[93]),
  .N7701(onet[94]),
  .N7702(onet[95]),
  .N7703(onet[96]),
  .N7704(onet[97]),
  .N7705(onet[98]),
  .N7706(onet[99]),
  .N7707(onet[100]),
  .N7735(onet[101]),
  .N7736(onet[102]),
  .N7737(onet[103]),
  .N7738(onet[104]),
  .N7739(onet[105]),
  .N7740(onet[106]),
  .N7741(onet[107]),
  .N7742(onet[108]),
  .N7754(onet[109]),
  .N7755(onet[110]),
  .N7756(onet[111]),
  .N7757(onet[112]),
  .N7758(onet[113]),
  .N7759(onet[114]),
  .N7760(onet[115]),
  .N7761(onet[116]),
  .N8075(onet[117]),
  .N8076(onet[118]),
  .N8123(onet[119]),
  .N8124(onet[120]),
  .N8127(onet[121]),
  .N8128(onet[122])
);

initial begin
  keepedCT = 0;
  totalCT = 0;
  uTests = 0; coverage = 0; 
  detectedFaultsAT =0; 
  faultIndex = 1; detectedListAT = 0; 
  expFCountCT = initialExpFCount; 
  testFile = $fopen("c5315-adj.tst", "w"); 
  #10; 

  while(coverage < desiredCoverage && uTests < utLimit) begin 
    detectedFaultsCT = 0; detectedListCT = 0;
    testVector = $random($time); 
    totalCT = totalCT + 1;
    uTests = uTests + 1; 
    faultIndex = 1; 
    #10; 
    newDiscovered = 0; 
    faultFile = $fopen ("c5315.flt", "r"); 
    while(!$feof(faultFile)) begin // Fault Injection loop 
      status=$fscanf(faultFile,"%s s@%b\n",wireName,stuckAtVal);  
      $InjectFault(wireName, stuckAtVal); 
      g = testVector;  
      #60;  
      
      if(o != onet) begin 
        detectedFaultsCT = detectedFaultsCT + 1;  
        detectedListCT[faultIndex] = 1'b1;  
        if(detectedListAT[faultIndex] == 0) begin 
          newDiscovered = newDiscovered + 1;
        end
      end //end of if 
      $RemoveFault(wireName); 
      #20;  
      faultIndex = faultIndex + 1;  
    end //end of while(!$feof(faultFile)) 
    $fclose(faultFile);
    
    if(newDiscovered < expFCountCT) begin
      tmp = expFCountCT / 2;
    end
    else begin
      tmp = (newDiscovered + expFCountCT) / 2; 
    end
    expFCountCT = tmp;  

    if(newDiscovered >= expFCountCT && (newDiscovered > 0)) begin 
      keepedCT = keepedCT + 1;
      uTests = 0;
      //detectedFaultsAT = 0; 
      detectedFaultsAT = detectedFaultsAT + newDiscovered; 
      for(faultIndex=1; faultIndex<=numOfFaults; faultIndex=faultIndex+1) 
        if(detectedListCT[faultIndex]==1) begin 
          $display ("here");
          detectedListAT[faultIndex] = 1'b1; 
        end 
             
      coverage = 100 * detectedFaultsAT / numOfFaults; 
      $fdisplay(testFile, "%b", testVector); 
    end
    #10; 
  end //end of while of Coverage 
	//	$display("Number of Random Vectors Generated: %d", uTests); 
  $display("%d of total %d test vectors are keeped!", keepedCT, totalCT);  
  $display("Coverage : %d", coverage); 
end

endmodule