`timescale 1ns / 1ps

module comparator (
  // Comparison Data
  input   logic [15:0]  Read_Data,
  input   logic [15:0]  Min_Reg,
  // Flags From Controller
  input   logic         Load_Min,
  // Flags To Min Registers
  output  logic         Load_Addr,
  output  logic         Load_Min_D
);

////////////////////////////////////////////////////////////////
///////////////////////   Internal Net   ///////////////////////
////////////////////////////////////////////////////////////////

logic lt;

////////////////////////////////////////////////////////////////
///////////////////////   Module Logic   ///////////////////////
////////////////////////////////////////////////////////////////

// Comparator
assign lt = (Read_Data < Min_Reg) ? 1'b1 : 1'b0;
assign Load_Min_D = (Load_Min | lt) ? 1'b1 : 1'b0;
assign Load_Addr = (Load_Min | lt) ? 1'b1 : 1'b0;

////////////////////////////////////////////////////////////////
//////////////////   Instantiation Template   //////////////////
////////////////////////////////////////////////////////////////
/*
comparator comparator (
  .Read_Data(),
  .Min_Reg(),
  .Load_Min(),
  .Load_Addr(),
  .Load_Min_D()
);
*/
endmodule