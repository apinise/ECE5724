
//Verilog file of module c5315
//CONVERTED BY CAD RESEARCH GROUP
//UNIVERSITY OF TEHRAN
//M. Hashem Haghbayan. hashem@cad.ut.ac.ir



`timescale 1 ns / 1ns

module c5315_net(

N1, 
N4, 
N11, 
N14, 
N17, 
N20, 
N23, 
N24, 
N25, 
N26, 
N27, 
N31, 
N34, 
N37, 
N40, 
N43, 
N46, 
N49, 
N52, 
N53, 
N54, 
N61, 
N64, 
N67, 
N70, 
N73, 
N76, 
N79, 
N80, 
N81, 
N82, 
N83, 
N86, 
N87, 
N88, 
N91, 
N94, 
N97, 
N100, 
N103, 
N106, 
N109, 
N112, 
N113, 
N114, 
N115, 
N116, 
N117, 
N118, 
N119, 
N120, 
N121, 
N122, 
N123, 
N126, 
N127, 
N128, 
N129, 
N130, 
N131, 
N132, 
N135, 
N136, 
N137, 
N140, 
N141, 
N145, 
N146, 
N149, 
N152, 
N155, 
N158, 
N161, 
N164, 
N167, 
N170, 
N173, 
N176, 
N179, 
N182, 
N185, 
N188, 
N191, 
N194, 
N197, 
N200, 
N203, 
N206, 
N209, 
N210, 
N217, 
N218, 
N225, 
N226, 
N233, 
N234, 
N241, 
N242, 
N245, 
N248, 
N251, 
N254, 
N257, 
N264, 
N265, 
N272, 
N273, 
N280, 
N281, 
N288, 
N289, 
N292, 
N293, 
N299, 
N302, 
N307, 
N308, 
N315, 
N316, 
N323, 
N324, 
N331, 
N332, 
N335, 
N338, 
N341, 
N348, 
N351, 
N358, 
N361, 
N366, 
N369, 
N372, 
N373, 
N374, 
N386, 
N389, 
N400, 
N411, 
N422, 
N435, 
N446, 
N457, 
N468, 
N479, 
N490, 
N503, 
N514, 
N523, 
N534, 
N545, 
N549, 
N552, 
N556, 
N559, 
N562, 
N566, 
N571, 
N574, 
N577, 
N580, 
N583, 
N588, 
N591, 
N592, 
N595, 
N596, 
N597, 
N598, 
N599, 
N603, 
N607, 
N610, 
N613, 
N616, 
N619, 
N625, 
N631, 

N709, 
N816, 
N1066, 
N1137, 
N1138, 
N1139, 
N1140, 
N1141, 
N1142, 
N1143, 
N1144, 
N1145, 
N1147, 
N1152, 
N1153, 
N1154, 
N1155, 
N1972, 
N2054, 
N2060, 
N2061, 
N2139, 
N2142, 
N2309, 
N2387, 
N2527, 
N2584, 
N2590, 
N2623, 
N3357, 
N3358, 
N3359, 
N3360, 
N3604, 
N3613, 
N4272, 
N4275, 
N4278, 
N4279, 
N4737, 
N4738, 
N4739, 
N4740, 
N5240, 
N5388, 
N6641, 
N6643, 
N6646, 
N6648, 
N6716, 
N6877, 
N6924, 
N6925, 
N6926, 
N6927, 
N7015, 
N7363, 
N7365, 
N7432, 
N7449, 
N7465, 
N7466, 
N7467, 
N7469, 
N7470, 
N7471, 
N7472, 
N7473, 
N7474, 
N7476, 
N7503, 
N7504, 
N7506, 
N7511, 
N7515, 
N7516, 
N7517, 
N7518, 
N7519, 
N7520, 
N7521, 
N7522, 
N7600, 
N7601, 
N7602, 
N7603, 
N7604, 
N7605, 
N7606, 
N7607, 
N7626, 
N7698, 
N7699, 
N7700, 
N7701, 
N7702, 
N7703, 
N7704, 
N7705, 
N7706, 
N7707, 
N7735, 
N7736, 
N7737, 
N7738, 
N7739, 
N7740, 
N7741, 
N7742, 
N7754, 
N7755, 
N7756, 
N7757, 
N7758, 
N7759, 
N7760, 
N7761, 
N8075, 
N8076, 
N8123, 
N8124, 
N8127, 
N8128);
input N1;
input N4;
input N11;
input N14;
input N17;
input N20;
input N23;
input N24;
input N25;
input N26;
input N27;
input N31;
input N34;
input N37;
input N40;
input N43;
input N46;
input N49;
input N52;
input N53;
input N54;
input N61;
input N64;
input N67;
input N70;
input N73;
input N76;
input N79;
input N80;
input N81;
input N82;
input N83;
input N86;
input N87;
input N88;
input N91;
input N94;
input N97;
input N100;
input N103;
input N106;
input N109;
input N112;
input N113;
input N114;
input N115;
input N116;
input N117;
input N118;
input N119;
input N120;
input N121;
input N122;
input N123;
input N126;
input N127;
input N128;
input N129;
input N130;
input N131;
input N132;
input N135;
input N136;
input N137;
input N140;
input N141;
input N145;
input N146;
input N149;
input N152;
input N155;
input N158;
input N161;
input N164;
input N167;
input N170;
input N173;
input N176;
input N179;
input N182;
input N185;
input N188;
input N191;
input N194;
input N197;
input N200;
input N203;
input N206;
input N209;
input N210;
input N217;
input N218;
input N225;
input N226;
input N233;
input N234;
input N241;
input N242;
input N245;
input N248;
input N251;
input N254;
input N257;
input N264;
input N265;
input N272;
input N273;
input N280;
input N281;
input N288;
input N289;
input N292;
input N293;
input N299;
input N302;
input N307;
input N308;
input N315;
input N316;
input N323;
input N324;
input N331;
input N332;
input N335;
input N338;
input N341;
input N348;
input N351;
input N358;
input N361;
input N366;
input N369;
input N372;
input N373;
input N374;
input N386;
input N389;
input N400;
input N411;
input N422;
input N435;
input N446;
input N457;
input N468;
input N479;
input N490;
input N503;
input N514;
input N523;
input N534;
input N545;
input N549;
input N552;
input N556;
input N559;
input N562;
input N566;
input N571;
input N574;
input N577;
input N580;
input N583;
input N588;
input N591;
input N592;
input N595;
input N596;
input N597;
input N598;
input N599;
input N603;
input N607;
input N610;
input N613;
input N616;
input N619;
input N625;
input N631;
output N709;
output N816;
output N1066;
output N1137;
output N1138;
output N1139;
output N1140;
output N1141;
output N1142;
output N1143;
output N1144;
output N1145;
output N1147;
output N1152;
output N1153;
output N1154;
output N1155;
output N1972;
output N2054;
output N2060;
output N2061;
output N2139;
output N2142;
output N2309;
output N2387;
output N2527;
output N2584;
output N2590;
output N2623;
output N3357;
output N3358;
output N3359;
output N3360;
output N3604;
output N3613;
output N4272;
output N4275;
output N4278;
output N4279;
output N4737;
output N4738;
output N4739;
output N4740;
output N5240;
output N5388;
output N6641;
output N6643;
output N6646;
output N6648;
output N6716;
output N6877;
output N6924;
output N6925;
output N6926;
output N6927;
output N7015;
output N7363;
output N7365;
output N7432;
output N7449;
output N7465;
output N7466;
output N7467;
output N7469;
output N7470;
output N7471;
output N7472;
output N7473;
output N7474;
output N7476;
output N7503;
output N7504;
output N7506;
output N7511;
output N7515;
output N7516;
output N7517;
output N7518;
output N7519;
output N7520;
output N7521;
output N7522;
output N7600;
output N7601;
output N7602;
output N7603;
output N7604;
output N7605;
output N7606;
output N7607;
output N7626;
output N7698;
output N7699;
output N7700;
output N7701;
output N7702;
output N7703;
output N7704;
output N7705;
output N7706;
output N7707;
output N7735;
output N7736;
output N7737;
output N7738;
output N7739;
output N7740;
output N7741;
output N7742;
output N7754;
output N7755;
output N7756;
output N7757;
output N7758;
output N7759;
output N7760;
output N7761;
output N8075;
output N8076;
output N8123;
output N8124;
output N8127;
output N8128;
wire
N1_0,
N1_1,
N4_0,
N4_1,
N4_2,
N4_3,
N4_4,
N4_5,
N11_0,
N11_1,
N14_0,
N14_1,
N17_0,
N17_1,
N20_0,
N20_1,
N27_0,
N27_1,
N27_2,
N31_0,
N31_1,
N34_0,
N34_1,
N37_0,
N37_1,
N40_0,
N40_1,
N43_0,
N43_1,
N46_0,
N46_1,
N49_0,
N49_1,
N54_0,
N54_1,
N54_2,
N54_3,
N54_4,
N54_5,
N61_0,
N61_1,
N64_0,
N64_1,
N67_0,
N67_1,
N70_0,
N70_1,
N73_0,
N73_1,
N76_0,
N76_1,
N83_0,
N83_1,
N88_0,
N88_1,
N91_0,
N91_1,
N94_0,
N94_1,
N97_0,
N97_1,
N100_0,
N100_1,
N103_0,
N103_1,
N106_0,
N106_1,
N109_0,
N109_1,
N123_0,
N123_1,
N132_0,
N132_1,
N137_0,
N137_1,
N141_0,
N141_1,
N141_2,
N146_0,
N146_1,
N149_0,
N149_1,
N152_0,
N152_1,
N155_0,
N155_1,
N158_0,
N158_1,
N161_0,
N161_1,
N164_0,
N164_1,
N167_0,
N167_1,
N170_0,
N170_1,
N173_0,
N173_1,
N176_0,
N176_1,
N179_0,
N179_1,
N182_0,
N182_1,
N185_0,
N185_1,
N188_0,
N188_1,
N191_0,
N191_1,
N194_0,
N194_1,
N197_0,
N197_1,
N200_0,
N200_1,
N203_0,
N203_1,
N206_0,
N206_1,
N210_0,
N210_1,
N210_2,
N210_3,
N210_4,
N210_5,
N218_0,
N218_1,
N218_2,
N218_3,
N218_4,
N218_5,
N226_0,
N226_1,
N226_2,
N226_3,
N226_4,
N226_5,
N234_0,
N234_1,
N234_2,
N234_3,
N234_4,
N234_5,
N242_0,
N242_1,
N245_0,
N245_1,
N248_0,
N248_1,
N251_0,
N251_1,
N254_0,
N254_1,
N257_0,
N257_1,
N257_2,
N257_3,
N257_4,
N257_5,
N265_0,
N265_1,
N265_2,
N265_3,
N265_4,
N265_5,
N273_0,
N273_1,
N273_2,
N273_3,
N273_4,
N273_5,
N281_0,
N281_1,
N281_2,
N281_3,
N281_4,
N281_5,
N289_0,
N289_1,
N293_0,
N293_1,
N293_2,
N293_3,
N293_4,
N299_0,
N299_1,
N302_0,
N302_1,
N302_2,
N302_3,
N308_0,
N308_1,
N308_2,
N308_3,
N308_4,
N308_5,
N316_0,
N316_1,
N316_2,
N316_3,
N316_4,
N316_5,
N324_0,
N324_1,
N324_2,
N324_3,
N324_4,
N324_5,
N332_0,
N332_1,
N335_0,
N335_1,
N338_0,
N338_1,
N341_0,
N341_1,
N341_2,
N341_3,
N341_4,
N341_5,
N348_0,
N348_1,
N351_0,
N351_1,
N351_2,
N351_3,
N351_4,
N351_5,
N358_0,
N358_1,
N361_0,
N361_1,
N361_2,
N361_3,
N366_0,
N366_1,
N369_0,
N369_1,
N374_0,
N374_1,
N374_2,
N374_3,
N374_4,
N374_5,
N374_6,
N374_7,
N374_8,
N374_9,
N374_10,
N386_0,
N386_1,
N389_0,
N389_1,
N389_2,
N389_3,
N389_4,
N389_5,
N389_6,
N389_7,
N389_8,
N389_9,
N400_0,
N400_1,
N400_2,
N400_3,
N400_4,
N400_5,
N400_6,
N400_7,
N400_8,
N400_9,
N411_0,
N411_1,
N411_2,
N411_3,
N411_4,
N411_5,
N411_6,
N411_7,
N411_8,
N411_9,
N422_0,
N422_1,
N422_2,
N422_3,
N422_4,
N422_5,
N422_6,
N422_7,
N422_8,
N422_9,
N422_10,
N422_11,
N435_0,
N435_1,
N435_2,
N435_3,
N435_4,
N435_5,
N435_6,
N435_7,
N435_8,
N435_9,
N446_0,
N446_1,
N446_2,
N446_3,
N446_4,
N446_5,
N446_6,
N446_7,
N446_8,
N446_9,
N457_0,
N457_1,
N457_2,
N457_3,
N457_4,
N457_5,
N457_6,
N457_7,
N457_8,
N457_9,
N468_0,
N468_1,
N468_2,
N468_3,
N468_4,
N468_5,
N468_6,
N468_7,
N468_8,
N468_9,
N479_0,
N479_1,
N479_2,
N479_3,
N479_4,
N479_5,
N479_6,
N479_7,
N479_8,
N479_9,
N490_0,
N490_1,
N490_2,
N490_3,
N490_4,
N490_5,
N490_6,
N490_7,
N490_8,
N490_9,
N490_10,
N490_11,
N503_0,
N503_1,
N503_2,
N503_3,
N503_4,
N503_5,
N503_6,
N503_7,
N503_8,
N503_9,
N514_0,
N514_1,
N514_2,
N514_3,
N514_4,
N514_5,
N514_6,
N514_7,
N523_0,
N523_1,
N523_2,
N523_3,
N523_4,
N523_5,
N523_6,
N523_7,
N523_8,
N523_9,
N534_0,
N534_1,
N534_2,
N534_3,
N534_4,
N534_5,
N534_6,
N534_7,
N534_8,
N534_9,
N545_0,
N545_1,
N545_2,
N549_0,
N549_1,
N552_0,
N552_1,
N552_2,
N556_0,
N556_1,
N559_0,
N559_1,
N562_0,
N562_1,
N562_2,
N566_0,
N566_1,
N566_2,
N566_3,
N571_0,
N571_1,
N574_0,
N574_1,
N577_0,
N577_1,
N580_0,
N580_1,
N583_0,
N583_1,
N583_2,
N583_3,
N588_0,
N588_1,
N592_0,
N592_1,
N599_0,
N599_1,
N599_2,
N603_0,
N603_1,
N603_2,
N607_0,
N607_1,
N610_0,
N610_1,
N613_0,
N613_1,
N616_0,
N616_1,
N619_0,
N619_1,
N619_2,
N619_3,
N619_4,
N625_0,
N625_1,
N625_2,
N625_3,
N625_4,
N1067_0,
N1067_1,
N1067_2,
N1067_3,
N1067_4,
N1067_5,
N1067_6,
N1067_7,
N1067_8,
N1067_9,
N1067_10,
N1067_11,
N1080_0,
N1080_1,
N1080_2,
N1080_3,
N1080_4,
N1080_5,
N1080_6,
N1080_7,
N1080_8,
N1080_9,
N1080_10,
N1092_0,
N1092_1,
N1092_2,
N1092_3,
N1092_4,
N1092_5,
N1092_6,
N1092_7,
N1092_8,
N1092_9,
N1092_10,
N1104_0,
N1104_1,
N1104_2,
N1104_3,
N1104_4,
N1104_5,
N1104_6,
N1104_7,
N1104_8,
N1104_9,
N1104_10,
N1104_11,
N1157_0,
N1157_1,
N1157_2,
N1161_0,
N1161_1,
N1161_2,
N1161_3,
N1161_4,
N1161_5,
N1161_6,
N1161_7,
N1161_8,
N1161_9,
N1161_10,
N1173_0,
N1173_1,
N1173_2,
N1173_3,
N1173_4,
N1173_5,
N1173_6,
N1173_7,
N1173_8,
N1173_9,
N1173_10,
N1185_0,
N1185_1,
N1185_2,
N1185_3,
N1185_4,
N1185_5,
N1185_6,
N1185_7,
N1185_8,
N1185_9,
N1185_10,
N1197_0,
N1197_1,
N1197_2,
N1197_3,
N1197_4,
N1197_5,
N1197_6,
N1197_7,
N1197_8,
N1197_9,
N1197_10,
N1209_0,
N1209_1,
N1209_2,
N1213_0,
N1213_1,
N1216_0,
N1216_1,
N1219_0,
N1219_1,
N1219_2,
N1223_0,
N1223_1,
N1223_2,
N1223_3,
N1223_4,
N1223_5,
N1223_6,
N1223_7,
N1223_8,
N1223_9,
N1223_10,
N1235_0,
N1235_1,
N1235_2,
N1235_3,
N1235_4,
N1235_5,
N1235_6,
N1235_7,
N1235_8,
N1235_9,
N1235_10,
N1247_0,
N1247_1,
N1247_2,
N1247_3,
N1247_4,
N1247_5,
N1247_6,
N1247_7,
N1247_8,
N1247_9,
N1247_10,
N1259_0,
N1259_1,
N1259_2,
N1259_3,
N1259_4,
N1259_5,
N1259_6,
N1259_7,
N1259_8,
N1259_9,
N1259_10,
N1271_0,
N1271_1,
N1271_2,
N1271_3,
N1271_4,
N1271_5,
N1271_6,
N1271_7,
N1280_0,
N1280_1,
N1280_2,
N1280_3,
N1280_4,
N1280_5,
N1280_6,
N1280_7,
N1280_8,
N1280_9,
N1280_10,
N1292_0,
N1292_1,
N1292_2,
N1292_3,
N1292_4,
N1292_5,
N1292_6,
N1292_7,
N1292_8,
N1292_9,
N1303_0,
N1303_1,
N1303_2,
N1303_3,
N1303_4,
N1303_5,
N1303_6,
N1303_7,
N1303_8,
N1303_9,
N1303_10,
N1315_0,
N1315_1,
N1315_2,
N1315_3,
N1315_4,
N1315_5,
N1315_6,
N1315_7,
N1315_8,
N1315_9,
N1315_10,
N1327_0,
N1327_1,
N1327_2,
N1327_3,
N1327_4,
N1327_5,
N1327_6,
N1327_7,
N1327_8,
N1327_9,
N1327_10,
N1339_0,
N1339_1,
N1339_2,
N1339_3,
N1339_4,
N1339_5,
N1339_6,
N1339_7,
N1339_8,
N1339_9,
N1339_10,
N1351_0,
N1351_1,
N1351_2,
N1351_3,
N1351_4,
N1351_5,
N1351_6,
N1351_7,
N1351_8,
N1351_9,
N1351_10,
N1363_0,
N1363_1,
N1363_2,
N1363_3,
N1363_4,
N1363_5,
N1363_6,
N1363_7,
N1363_8,
N1363_9,
N1363_10,
N1375_0,
N1375_1,
N1378_0,
N1378_1,
N1381_0,
N1381_1,
N1384_0,
N1384_1,
N1387_0,
N1387_1,
N1390_0,
N1390_1,
N1393_0,
N1393_1,
N1396_0,
N1396_1,
N1415_0,
N1415_1,
N1418_0,
N1418_1,
N1421_0,
N1421_1,
N1424_0,
N1424_1,
N1427_0,
N1427_1,
N1430_0,
N1430_1,
N1433_0,
N1433_1,
N1436_0,
N1436_1,
N1455_0,
N1455_1,
N1455_2,
N1455_3,
N1455_4,
N1455_5,
N1462_0,
N1462_1,
N1462_2,
N1462_3,
N1462_4,
N1462_5,
N1469_0,
N1469_1,
N1469_2,
N1469_3,
N1469_4,
N1475_0,
N1475_1,
N1475_2,
N1479_0,
N1479_1,
N1482_0,
N1482_1,
N1482_2,
N1482_3,
N1482_4,
N1482_5,
N1482_6,
N1482_7,
N1482_8,
N1492_0,
N1492_1,
N1495_0,
N1495_1,
N1498_0,
N1498_1,
N1501_0,
N1501_1,
N1504_0,
N1504_1,
N1507_0,
N1507_1,
N1510_0,
N1510_1,
N1513_0,
N1513_1,
N1516_0,
N1516_1,
N1519_0,
N1519_1,
N1522_0,
N1522_1,
N1525_0,
N1525_1,
N1542_0,
N1542_1,
N1545_0,
N1545_1,
N1548_0,
N1548_1,
N1551_0,
N1551_1,
N1554_0,
N1554_1,
N1557_0,
N1557_1,
N1560_0,
N1560_1,
N1563_0,
N1563_1,
N1566_0,
N1566_1,
N1566_2,
N1566_3,
N1566_4,
N1566_5,
N1573_0,
N1573_1,
N1573_2,
N1573_3,
N1573_4,
N1573_5,
N1580_0,
N1580_1,
N1583_0,
N1583_1,
N1583_2,
N1583_3,
N1588_0,
N1588_1,
N1588_2,
N1588_3,
N1588_4,
N1594_0,
N1594_1,
N1597_0,
N1597_1,
N1600_0,
N1600_1,
N1603_0,
N1603_1,
N1606_0,
N1606_1,
N1609_0,
N1609_1,
N1612_0,
N1612_1,
N1615_0,
N1615_1,
N1618_0,
N1618_1,
N1621_0,
N1621_1,
N1624_0,
N1624_1,
N1627_0,
N1627_1,
N1630_0,
N1630_1,
N1633_0,
N1633_1,
N1636_0,
N1636_1,
N1639_0,
N1639_1,
N1642_0,
N1642_1,
N1645_0,
N1645_1,
N1648_0,
N1648_1,
N1651_0,
N1651_1,
N1654_0,
N1654_1,
N1657_0,
N1657_1,
N1660_0,
N1660_1,
N1663_0,
N1663_1,
N1663_2,
N1663_3,
N1663_4,
N1663_5,
N1663_6,
N1663_7,
N1663_8,
N1663_9,
N1663_10,
N1675_0,
N1675_1,
N1675_2,
N1675_3,
N1675_4,
N1675_5,
N1675_6,
N1675_7,
N1675_8,
N1685_0,
N1685_1,
N1685_2,
N1685_3,
N1685_4,
N1685_5,
N1685_6,
N1685_7,
N1685_8,
N1685_9,
N1685_10,
N1697_0,
N1697_1,
N1697_2,
N1697_3,
N1697_4,
N1697_5,
N1697_6,
N1697_7,
N1697_8,
N1697_9,
N1697_10,
N1709_0,
N1709_1,
N1709_2,
N1709_3,
N1709_4,
N1709_5,
N1709_6,
N1709_7,
N1709_8,
N1709_9,
N1709_10,
N1721_0,
N1721_1,
N1721_2,
N1721_3,
N1721_4,
N1727_0,
N1727_1,
N1727_2,
N1731_0,
N1731_1,
N1731_2,
N1731_3,
N1731_4,
N1731_5,
N1731_6,
N1731_7,
N1731_8,
N1731_9,
N1731_10,
N1743_0,
N1743_1,
N1743_2,
N1743_3,
N1743_4,
N1743_5,
N1743_6,
N1743_7,
N1743_8,
N1743_9,
N1743_10,
N1755_0,
N1755_1,
N1758_0,
N1758_1,
N1761_0,
N1761_1,
N1761_2,
N1761_3,
N1761_4,
N1761_5,
N1761_6,
N1769_0,
N1769_1,
N1769_2,
N1769_3,
N1769_4,
N1769_5,
N1769_6,
N1777_0,
N1777_1,
N1777_2,
N1777_3,
N1777_4,
N1777_5,
N1777_6,
N1785_0,
N1785_1,
N1785_2,
N1785_3,
N1785_4,
N1785_5,
N1785_6,
N1793_0,
N1793_1,
N1793_2,
N1793_3,
N1793_4,
N1793_5,
N1800_0,
N1800_1,
N1800_2,
N1800_3,
N1800_4,
N1800_5,
N1807_0,
N1807_1,
N1807_2,
N1807_3,
N1807_4,
N1807_5,
N1814_0,
N1814_1,
N1814_2,
N1814_3,
N1814_4,
N1814_5,
N1821_0,
N1821_1,
N1824_0,
N1824_1,
N1827_0,
N1827_1,
N1830_0,
N1830_1,
N1833_0,
N1833_1,
N1836_0,
N1836_1,
N1839_0,
N1839_1,
N1842_0,
N1842_1,
N1845_0,
N1845_1,
N1848_0,
N1848_1,
N1851_0,
N1851_1,
N1854_0,
N1854_1,
N1857_0,
N1857_1,
N1860_0,
N1860_1,
N1863_0,
N1863_1,
N1866_0,
N1866_1,
N1869_0,
N1869_1,
N1872_0,
N1872_1,
N1875_0,
N1875_1,
N1878_0,
N1878_1,
N1881_0,
N1881_1,
N1884_0,
N1884_1,
N1887_0,
N1887_1,
N1890_0,
N1890_1,
N1893_0,
N1893_1,
N1896_0,
N1896_1,
N1899_0,
N1899_1,
N1902_0,
N1902_1,
N1905_0,
N1905_1,
N1908_0,
N1908_1,
N1911_0,
N1911_1,
N1914_0,
N1914_1,
N1917_0,
N1917_1,
N1920_0,
N1920_1,
N1923_0,
N1923_1,
N1926_0,
N1926_1,
N1929_0,
N1929_1,
N1932_0,
N1932_1,
N1935_0,
N1935_1,
N1938_0,
N1938_1,
N1941_0,
N1941_1,
N1944_0,
N1944_1,
N1947_0,
N1947_1,
N1950_0,
N1950_1,
N1953_0,
N1953_1,
N1956_0,
N1956_1,
N1959_0,
N1959_1,
N1962_0,
N1962_1,
N1965_0,
N1965_1,
N1968_0,
N1968_1,
N2647_0,
N2647_1,
N2647_2,
N2647_3,
N2647_4,
N2653_0,
N2653_1,
N2653_2,
N2653_3,
N2653_4,
N2653_5,
N2653_6,
N2653_7,
N2653_8,
N2653_9,
N2664_0,
N2664_1,
N2664_2,
N2664_3,
N2664_4,
N2664_5,
N2664_6,
N2664_7,
N2664_8,
N2664_9,
N2675_0,
N2675_1,
N2675_2,
N2675_3,
N2675_4,
N2681_0,
N2681_1,
N2681_2,
N2681_3,
N2681_4,
N2681_5,
N2681_6,
N2681_7,
N2681_8,
N2681_9,
N2692_0,
N2692_1,
N2692_2,
N2692_3,
N2692_4,
N2692_5,
N2692_6,
N2692_7,
N2692_8,
N2692_9,
N2704_0,
N2704_1,
N2704_2,
N2704_3,
N2722_0,
N2722_1,
N2722_2,
N2722_3,
N2722_4,
N2728_0,
N2728_1,
N2728_2,
N2728_3,
N2728_4,
N2728_5,
N2728_6,
N2728_7,
N2728_8,
N2728_9,
N2739_0,
N2739_1,
N2739_2,
N2739_3,
N2739_4,
N2739_5,
N2739_6,
N2739_7,
N2739_8,
N2739_9,
N2750_0,
N2750_1,
N2750_2,
N2750_3,
N2750_4,
N2756_0,
N2756_1,
N2756_2,
N2756_3,
N2756_4,
N2756_5,
N2756_6,
N2756_7,
N2756_8,
N2756_9,
N2767_0,
N2767_1,
N2767_2,
N2767_3,
N2767_4,
N2767_5,
N2767_6,
N2767_7,
N2767_8,
N2767_9,
N2779_0,
N2779_1,
N2779_2,
N2779_3,
N2779_4,
N2779_5,
N2779_6,
N2779_7,
N2779_8,
N2779_9,
N2790_0,
N2790_1,
N2790_2,
N2790_3,
N2790_4,
N2790_5,
N2790_6,
N2790_7,
N2790_8,
N2790_9,
N2801_0,
N2801_1,
N2801_2,
N2801_3,
N2801_4,
N2801_5,
N2801_6,
N2801_7,
N2801_8,
N2801_9,
N2812_0,
N2812_1,
N2812_2,
N2812_3,
N2812_4,
N2812_5,
N2812_6,
N2812_7,
N2812_8,
N2812_9,
N2855_0,
N2855_1,
N2855_2,
N2855_3,
N2855_4,
N2861_0,
N2861_1,
N2861_2,
N2861_3,
N2861_4,
N2877_0,
N2877_1,
N2877_2,
N2877_3,
N2882_0,
N2882_1,
N2882_2,
N2882_3,
N2882_4,
N2882_5,
N2882_6,
N2882_7,
N2891_0,
N2891_1,
N2891_2,
N2891_3,
N2891_4,
N2891_5,
N2891_6,
N2891_7,
N2891_8,
N2942_0,
N2942_1,
N2942_2,
N2942_3,
N2942_4,
N2948_0,
N2948_1,
N2948_2,
N2948_3,
N2948_4,
N2964_0,
N2964_1,
N2964_2,
N2964_3,
N3000_0,
N3000_1,
N3003_0,
N3003_1,
N3007_0,
N3007_1,
N3010_0,
N3010_1,
N3035_0,
N3035_1,
N3038_0,
N3038_1,
N3041_0,
N3041_1,
N3041_2,
N3041_3,
N3041_4,
N3041_5,
N3041_6,
N3041_7,
N3041_8,
N3041_9,
N3052_0,
N3052_1,
N3052_2,
N3052_3,
N3052_4,
N3052_5,
N3052_6,
N3052_7,
N3052_8,
N3052_9,
N3063_0,
N3063_1,
N3063_2,
N3063_3,
N3068_0,
N3068_1,
N3075_0,
N3075_1,
N3075_2,
N3075_3,
N3075_4,
N3075_5,
N3075_6,
N3075_7,
N3075_8,
N3075_9,
N3086_0,
N3086_1,
N3086_2,
N3086_3,
N3086_4,
N3086_5,
N3086_6,
N3086_7,
N3086_8,
N3086_9,
N3097_0,
N3097_1,
N3097_2,
N3097_3,
N3097_4,
N3097_5,
N3097_6,
N3097_7,
N3097_8,
N3097_9,
N3108_0,
N3108_1,
N3108_2,
N3108_3,
N3108_4,
N3108_5,
N3108_6,
N3108_7,
N3108_8,
N3108_9,
N3119_0,
N3119_1,
N3119_2,
N3119_3,
N3119_4,
N3119_5,
N3119_6,
N3119_7,
N3119_8,
N3119_9,
N3130_0,
N3130_1,
N3130_2,
N3130_3,
N3130_4,
N3130_5,
N3130_6,
N3130_7,
N3130_8,
N3130_9,
N3147_0,
N3147_1,
N3147_2,
N3147_3,
N3147_4,
N3147_5,
N3147_6,
N3147_7,
N3147_8,
N3147_9,
N3158_0,
N3158_1,
N3158_2,
N3158_3,
N3158_4,
N3158_5,
N3158_6,
N3158_7,
N3158_8,
N3158_9,
N3169_0,
N3169_1,
N3169_2,
N3169_3,
N3169_4,
N3169_5,
N3169_6,
N3169_7,
N3169_8,
N3169_9,
N3180_0,
N3180_1,
N3180_2,
N3180_3,
N3180_4,
N3180_5,
N3180_6,
N3180_7,
N3180_8,
N3180_9,
N3191_0,
N3191_1,
N3200_0,
N3200_1,
N3456_0,
N3456_1,
N3691_0,
N3691_1,
N3691_2,
N3691_3,
N3691_4,
N3691_5,
N3691_6,
N3691_7,
N3705_0,
N3705_1,
N3732_0,
N3732_1,
N3732_2,
N3732_3,
N3732_4,
N3771_0,
N3771_1,
N3771_2,
N3775_0,
N3775_1,
N3775_2,
N3789_0,
N3789_1,
N3789_2,
N3793_0,
N3793_1,
N3793_2,
N3797_0,
N3797_1,
N3810_0,
N3810_1,
N3813_0,
N3813_1,
N3816_0,
N3816_1,
N3819_0,
N3819_1,
N3824_0,
N3824_1,
N3842_0,
N3842_1,
N3842_2,
N3842_3,
N3842_4,
N3842_5,
N3849_0,
N3849_1,
N3849_2,
N3849_3,
N3849_4,
N3855_0,
N3855_1,
N3855_2,
N3855_3,
N3855_4,
N3861_0,
N3861_1,
N3861_2,
N3861_3,
N3861_4,
N3867_0,
N3867_1,
N3867_2,
N3867_3,
N3867_4,
N3873_0,
N3873_1,
N3873_2,
N3873_3,
N3873_4,
N3873_5,
N3873_6,
N3881_0,
N3881_1,
N3881_2,
N3881_3,
N3881_4,
N3887_0,
N3887_1,
N3887_2,
N3887_3,
N3887_4,
N3893_0,
N3893_1,
N3893_2,
N3893_3,
N3893_4,
N3911_0,
N3911_1,
N3921_0,
N3921_1,
N3921_2,
N3921_3,
N3921_4,
N3927_0,
N3927_1,
N3927_2,
N3927_3,
N3927_4,
N3933_0,
N3933_1,
N3933_2,
N3933_3,
N3933_4,
N3942_0,
N3942_1,
N3942_2,
N3942_3,
N3942_4,
N3948_0,
N3948_1,
N3948_2,
N3948_3,
N3948_4,
N3948_5,
N3948_6,
N3956_0,
N3956_1,
N3956_2,
N3956_3,
N3956_4,
N3962_0,
N3962_1,
N3962_2,
N3962_3,
N3962_4,
N3968_0,
N3968_1,
N3968_2,
N3968_3,
N3968_4,
N3968_5,
N3984_0,
N3984_1,
N4008_0,
N4008_1,
N4011_0,
N4011_1,
N4021_0,
N4021_1,
N4067_0,
N4067_1,
N4080_0,
N4080_1,
N4080_2,
N4088_0,
N4088_1,
N4091_0,
N4091_1,
N4094_0,
N4094_1,
N4097_0,
N4097_1,
N4100_0,
N4100_1,
N4103_0,
N4103_1,
N4106_0,
N4106_1,
N4109_0,
N4109_1,
N4144_0,
N4144_1,
N4147_0,
N4147_1,
N4150_0,
N4150_1,
N4153_0,
N4153_1,
N4156_0,
N4156_1,
N4159_0,
N4159_1,
N4188_0,
N4188_1,
N4191_0,
N4191_1,
N4200_0,
N4200_1,
N4203_0,
N4203_1,
N4206_0,
N4206_1,
N4209_0,
N4209_1,
N4212_0,
N4212_1,
N4215_0,
N4215_1,
N4219_0,
N4219_1,
N4225_0,
N4225_1,
N4228_0,
N4228_1,
N4231_0,
N4231_1,
N4234_0,
N4234_1,
N4237_0,
N4237_1,
N4240_0,
N4240_1,
N4243_0,
N4243_1,
N4246_0,
N4246_1,
N4249_0,
N4249_1,
N4252_0,
N4252_1,
N4255_0,
N4255_1,
N4258_0,
N4258_1,
N4264_0,
N4264_1,
N4280_0,
N4280_1,
N4280_2,
N4284_0,
N4284_1,
N4284_2,
N4284_3,
N4284_4,
N4290_0,
N4290_1,
N4290_2,
N4290_3,
N4290_4,
N4290_5,
N4298_0,
N4298_1,
N4301_0,
N4301_1,
N4301_2,
N4305_0,
N4305_1,
N4305_2,
N4305_3,
N4310_0,
N4310_1,
N4310_2,
N4310_3,
N4310_4,
N4316_0,
N4316_1,
N4316_2,
N4320_0,
N4320_1,
N4320_2,
N4320_3,
N4325_0,
N4325_1,
N4325_2,
N4325_3,
N4325_4,
N4332_0,
N4332_1,
N4332_2,
N4336_0,
N4336_1,
N4336_2,
N4336_3,
N4336_4,
N4342_0,
N4342_1,
N4342_2,
N4342_3,
N4342_4,
N4342_5,
N4349_0,
N4349_1,
N4349_2,
N4349_3,
N4349_4,
N4349_5,
N4349_6,
N4357_0,
N4357_1,
N4357_2,
N4357_3,
N4357_4,
N4357_5,
N4364_0,
N4364_1,
N4364_2,
N4364_3,
N4364_4,
N4364_5,
N4364_6,
N4364_7,
N4364_8,
N4364_9,
N4375_0,
N4375_1,
N4375_2,
N4379_0,
N4379_1,
N4379_2,
N4379_3,
N4379_4,
N4385_0,
N4385_1,
N4385_2,
N4385_3,
N4385_4,
N4385_5,
N4396_0,
N4396_1,
N4396_2,
N4400_0,
N4400_1,
N4400_2,
N4400_3,
N4405_0,
N4405_1,
N4405_2,
N4405_3,
N4405_4,
N4405_5,
N4412_0,
N4412_1,
N4412_2,
N4412_3,
N4412_4,
N4418_0,
N4418_1,
N4418_2,
N4418_3,
N4418_4,
N4418_5,
N4425_0,
N4425_1,
N4425_2,
N4425_3,
N4425_4,
N4425_5,
N4425_6,
N4425_7,
N4425_8,
N4425_9,
N4436_0,
N4436_1,
N4436_2,
N4440_0,
N4440_1,
N4440_2,
N4440_3,
N4445_0,
N4445_1,
N4445_2,
N4445_3,
N4445_4,
N4456_0,
N4456_1,
N4456_2,
N4456_3,
N4456_4,
N4462_0,
N4462_1,
N4462_2,
N4462_3,
N4462_4,
N4462_5,
N4469_0,
N4469_1,
N4469_2,
N4469_3,
N4469_4,
N4469_5,
N4469_6,
N4477_0,
N4477_1,
N4477_2,
N4477_3,
N4477_4,
N4477_5,
N4512_0,
N4512_1,
N4524_0,
N4524_1,
N4524_2,
N4532_0,
N4532_1,
N4532_2,
N4548_0,
N4548_1,
N4551_0,
N4551_1,
N4554_0,
N4554_1,
N4557_0,
N4557_1,
N4560_0,
N4560_1,
N4563_0,
N4563_1,
N4566_0,
N4566_1,
N4569_0,
N4569_1,
N4572_0,
N4572_1,
N4575_0,
N4575_1,
N4578_0,
N4578_1,
N4581_0,
N4581_1,
N4584_0,
N4584_1,
N4587_0,
N4587_1,
N4590_0,
N4590_1,
N4593_0,
N4593_1,
N4596_0,
N4596_1,
N4599_0,
N4599_1,
N4602_0,
N4602_1,
N4605_0,
N4605_1,
N4608_0,
N4608_1,
N4611_0,
N4611_1,
N4614_0,
N4614_1,
N4617_0,
N4617_1,
N4621_0,
N4621_1,
N4624_0,
N4624_1,
N4627_0,
N4627_1,
N4630_0,
N4630_1,
N4633_0,
N4633_1,
N4637_0,
N4637_1,
N4640_0,
N4640_1,
N4643_0,
N4643_1,
N4646_0,
N4646_1,
N4649_0,
N4649_1,
N4652_0,
N4652_1,
N4655_0,
N4655_1,
N4658_0,
N4658_1,
N4662_0,
N4662_1,
N4665_0,
N4665_1,
N4668_0,
N4668_1,
N4671_0,
N4671_1,
N4674_0,
N4674_1,
N4677_0,
N4677_1,
N4680_0,
N4680_1,
N4683_0,
N4683_1,
N4686_0,
N4686_1,
N4689_0,
N4689_1,
N4692_0,
N4692_1,
N4695_0,
N4695_1,
N4698_0,
N4698_1,
N4939_0,
N4939_1,
N5049_0,
N5049_1,
N5150_0,
N5150_1,
N5157_0,
N5157_1,
N5166_0,
N5166_1,
N5169_0,
N5169_1,
N5173_0,
N5173_1,
N5177_0,
N5177_1,
N5180_0,
N5180_1,
N5183_0,
N5183_1,
N5186_0,
N5186_1,
N5189_0,
N5189_1,
N5192_0,
N5192_1,
N5195_0,
N5195_1,
N5199_0,
N5199_1,
N5202_0,
N5202_1,
N5205_0,
N5205_1,
N5208_0,
N5208_1,
N5211_0,
N5211_1,
N5214_0,
N5214_1,
N5217_0,
N5217_1,
N5220_0,
N5220_1,
N5236_0,
N5236_1,
N5264_0,
N5264_1,
N5264_2,
N5264_3,
N5264_4,
N5264_5,
N5264_6,
N5264_7,
N5264_8,
N5284_0,
N5284_1,
N5284_2,
N5284_3,
N5284_4,
N5284_5,
N5284_6,
N5284_7,
N5284_8,
N5284_9,
N5284_10,
N5284_11,
N5284_12,
N5315_0,
N5315_1,
N5315_2,
N5319_0,
N5319_1,
N5324_0,
N5324_1,
N5324_2,
N5328_0,
N5328_1,
N5346_0,
N5346_1,
N5371_0,
N5371_1,
N5374_0,
N5374_1,
N5377_0,
N5377_1,
N5382_0,
N5382_1,
N5385_0,
N5385_1,
N5389_0,
N5389_1,
N5389_2,
N5389_3,
N5389_4,
N5389_5,
N5396_0,
N5396_1,
N5396_2,
N5396_3,
N5396_4,
N5396_5,
N5396_6,
N5396_7,
N5396_8,
N5396_9,
N5407_0,
N5407_1,
N5407_2,
N5407_3,
N5407_4,
N5407_5,
N5407_6,
N5407_7,
N5407_8,
N5407_9,
N5418_0,
N5418_1,
N5418_2,
N5418_3,
N5418_4,
N5424_0,
N5424_1,
N5424_2,
N5424_3,
N5424_4,
N5424_5,
N5431_0,
N5431_1,
N5431_2,
N5431_3,
N5431_4,
N5431_5,
N5431_6,
N5431_7,
N5431_8,
N5441_0,
N5441_1,
N5441_2,
N5441_3,
N5441_4,
N5441_5,
N5441_6,
N5441_7,
N5441_8,
N5441_9,
N5452_0,
N5452_1,
N5452_2,
N5452_3,
N5452_4,
N5452_5,
N5452_6,
N5452_7,
N5452_8,
N5462_0,
N5462_1,
N5462_2,
N5462_3,
N5462_4,
N5462_5,
N5470_0,
N5470_1,
N5470_2,
N5470_3,
N5470_4,
N5470_5,
N5477_0,
N5477_1,
N5477_2,
N5477_3,
N5477_4,
N5477_5,
N5477_6,
N5477_7,
N5477_8,
N5477_9,
N5488_0,
N5488_1,
N5488_2,
N5488_3,
N5488_4,
N5488_5,
N5488_6,
N5488_7,
N5488_8,
N5498_0,
N5498_1,
N5498_2,
N5498_3,
N5498_4,
N5498_5,
N5498_6,
N5506_0,
N5506_1,
N5506_2,
N5506_3,
N5506_4,
N5506_5,
N5506_6,
N5506_7,
N5506_8,
N5506_9,
N5506_10,
N5506_11,
N5506_12,
N5520_0,
N5520_1,
N5520_2,
N5520_3,
N5520_4,
N5520_5,
N5520_6,
N5520_7,
N5520_8,
N5520_9,
N5520_10,
N5520_11,
N5520_12,
N5520_13,
N5520_14,
N5536_0,
N5536_1,
N5536_2,
N5536_3,
N5536_4,
N5536_5,
N5536_6,
N5536_7,
N5536_8,
N5536_9,
N5536_10,
N5536_11,
N5549_0,
N5549_1,
N5549_2,
N5549_3,
N5549_4,
N5555_0,
N5555_1,
N5555_2,
N5555_3,
N5555_4,
N5555_5,
N5562_0,
N5562_1,
N5562_2,
N5562_3,
N5562_4,
N5562_5,
N5562_6,
N5562_7,
N5562_8,
N5562_9,
N5573_0,
N5573_1,
N5573_2,
N5573_3,
N5573_4,
N5579_0,
N5579_1,
N5579_2,
N5579_3,
N5579_4,
N5579_5,
N5595_0,
N5595_1,
N5595_2,
N5595_3,
N5595_4,
N5595_5,
N5595_6,
N5595_7,
N5595_8,
N5595_9,
N5606_0,
N5606_1,
N5606_2,
N5606_3,
N5606_4,
N5606_5,
N5606_6,
N5606_7,
N5606_8,
N5624_0,
N5624_1,
N5624_2,
N5624_3,
N5624_4,
N5624_5,
N5624_6,
N5624_7,
N5624_8,
N5634_0,
N5634_1,
N5634_2,
N5634_3,
N5634_4,
N5634_5,
N5634_6,
N5655_0,
N5655_1,
N5655_2,
N5655_3,
N5655_4,
N5655_5,
N5655_6,
N5655_7,
N5655_8,
N5655_9,
N5655_10,
N5655_11,
N5655_12,
N5655_13,
N5655_14,
N5671_0,
N5671_1,
N5671_2,
N5671_3,
N5671_4,
N5671_5,
N5671_6,
N5671_7,
N5671_8,
N5671_9,
N5671_10,
N5671_11,
N5684_0,
N5684_1,
N5684_2,
N5684_3,
N5684_4,
N5692_0,
N5692_1,
N5692_2,
N5696_0,
N5696_1,
N5696_2,
N5700_0,
N5700_1,
N5703_0,
N5703_1,
N5703_2,
N5707_0,
N5707_1,
N5707_2,
N5711_0,
N5711_1,
N5736_0,
N5736_1,
N5739_0,
N5739_1,
N5742_0,
N5742_1,
N5745_0,
N5745_1,
N5756_0,
N5756_1,
N6025_0,
N6025_1,
N6028_0,
N6028_1,
N6031_0,
N6031_1,
N6034_0,
N6034_1,
N6037_0,
N6037_1,
N6040_0,
N6040_1,
N6045_0,
N6045_1,
N6048_0,
N6048_1,
N6051_0,
N6051_1,
N6054_0,
N6054_1,
N6080_0,
N6080_1,
N6091_0,
N6091_1,
N6108_0,
N6108_1,
N6117_0,
N6117_1,
N6140_0,
N6140_1,
N6149_0,
N6149_1,
N6164_0,
N6164_1,
N6168_0,
N6168_1,
N6175_0,
N6175_1,
N6197_0,
N6197_1,
N6200_0,
N6200_1,
N6203_0,
N6203_1,
N6206_0,
N6206_1,
N6209_0,
N6209_1,
N6212_0,
N6212_1,
N6215_0,
N6215_1,
N6218_0,
N6218_1,
N6238_0,
N6238_1,
N6241_0,
N6241_1,
N6244_0,
N6244_1,
N6247_0,
N6247_1,
N6250_0,
N6250_1,
N6253_0,
N6253_1,
N6256_0,
N6256_1,
N6259_0,
N6259_1,
N6262_0,
N6262_1,
N6265_0,
N6265_1,
N6268_0,
N6268_1,
N6271_0,
N6271_1,
N6274_0,
N6274_1,
N6277_0,
N6277_1,
N6280_0,
N6280_1,
N6283_0,
N6283_1,
N6286_0,
N6286_1,
N6289_0,
N6289_1,
N6292_0,
N6292_1,
N6295_0,
N6295_1,
N6298_0,
N6298_1,
N6301_0,
N6301_1,
N6304_0,
N6304_1,
N6307_0,
N6307_1,
N6310_0,
N6310_1,
N6313_0,
N6313_1,
N6316_0,
N6316_1,
N6319_0,
N6319_1,
N6322_0,
N6322_1,
N6325_0,
N6325_1,
N6328_0,
N6328_1,
N6331_0,
N6331_1,
N6335_0,
N6335_1,
N6338_0,
N6338_1,
N6341_0,
N6341_1,
N6344_0,
N6344_1,
N6347_0,
N6347_1,
N6350_0,
N6350_1,
N6353_0,
N6353_1,
N6356_0,
N6356_1,
N6359_0,
N6359_1,
N6364_0,
N6364_1,
N6367_0,
N6367_1,
N6370_0,
N6370_1,
N6397_0,
N6397_1,
N6411_0,
N6411_1,
N6415_0,
N6415_1,
N6415_2,
N6419_0,
N6419_1,
N6427_0,
N6427_1,
N6437_0,
N6437_1,
N6441_0,
N6441_1,
N6441_2,
N6445_0,
N6445_1,
N6466_0,
N6466_1,
N6478_0,
N6478_1,
N6482_0,
N6482_1,
N6486_0,
N6486_1,
N6490_0,
N6490_1,
N6494_0,
N6494_1,
N6500_0,
N6500_1,
N6504_0,
N6504_1,
N6508_0,
N6508_1,
N6512_0,
N6512_1,
N6516_0,
N6516_1,
N6526_0,
N6526_1,
N6536_0,
N6536_1,
N6539_0,
N6539_1,
N6553_0,
N6553_1,
N6556_0,
N6556_1,
N6566_0,
N6566_1,
N6569_0,
N6569_1,
N6572_0,
N6572_1,
N6575_0,
N6575_1,
N6580_0,
N6580_1,
N6584_0,
N6584_1,
N6587_0,
N6587_1,
N6592_0,
N6592_1,
N6599_0,
N6599_1,
N6606_0,
N6606_1,
N6609_0,
N6609_1,
N6619_0,
N6619_1,
N6622_0,
N6622_1,
N6634_0,
N6634_1,
N6637_0,
N6637_1,
N6724_0,
N6724_1,
N6792_0,
N6792_1,
N6795_0,
N6795_1,
N6817_0,
N6817_1,
N6817_2,
N6817_3,
N6817_4,
N6831_0,
N6831_1,
N6844_0,
N6844_1,
N6844_2,
N6844_3,
N6844_4,
N6857_0,
N6857_1,
N6866_0,
N6866_1,
N6866_2,
N6866_3,
N6866_4,
N6881_0,
N6881_1,
N6885_0,
N6885_1,
N6891_0,
N6891_1,
N6897_0,
N6897_1,
N6901_0,
N6901_1,
N6905_0,
N6905_1,
N6909_0,
N6909_1,
N6916_0,
N6916_1,
N6932_0,
N6932_1,
N6967_0,
N6967_1,
N6979_0,
N6979_1,
N6979_2,
N7003_0,
N7003_1,
N7006_0,
N7006_1,
N7023_0,
N7023_1,
N7023_2,
N7023_3,
N7028_0,
N7028_1,
N7031_0,
N7031_1,
N7034_0,
N7034_1,
N7037_0,
N7037_1,
N7041_0,
N7041_1,
N7049_0,
N7049_1,
N7049_2,
N7049_3,
N7054_0,
N7054_1,
N7057_0,
N7057_1,
N7060_0,
N7060_1,
N7065_0,
N7065_1,
N7076_0,
N7076_1,
N7080_0,
N7080_1,
N7090_0,
N7090_1,
N7094_0,
N7094_1,
N7097_0,
N7097_1,
N7101_0,
N7101_1,
N7190_0,
N7190_1,
N7190_2,
N7190_3,
N7190_4,
N7198_0,
N7198_1,
N7198_2,
N7198_3,
N7198_4,
N7209_0,
N7209_1,
N7212_0,
N7212_1,
N7219_0,
N7219_1,
N7222_0,
N7222_1,
N7225_0,
N7225_1,
N7236_0,
N7236_1,
N7239_0,
N7239_1,
N7242_0,
N7242_1,
N7245_0,
N7245_1,
N7250_0,
N7250_1,
N7250_2,
N7250_3,
N7250_4,
N7250_5,
N7257_0,
N7257_1,
N7260_0,
N7260_1,
N7263_0,
N7263_1,
N7270_0,
N7270_1,
N7270_2,
N7270_3,
N7270_4,
N7276_0,
N7276_1,
N7276_2,
N7276_3,
N7276_4,
N7282_0,
N7282_1,
N7282_2,
N7282_3,
N7282_4,
N7288_0,
N7288_1,
N7288_2,
N7288_3,
N7288_4,
N7294_0,
N7294_1,
N7294_2,
N7294_3,
N7294_4,
N7301_0,
N7301_1,
N7304_0,
N7304_1,
N7304_2,
N7304_3,
N7304_4,
N7310_0,
N7310_1,
N7310_2,
N7310_3,
N7310_4,
N7394_0,
N7394_1,
N7397_0,
N7397_1,
N7402_0,
N7402_1,
N7409_0,
N7409_1,
N7412_0,
N7412_1,
N7421_0,
N7421_1,
N7489_0,
N7489_1,
N7531_0,
N7531_1,
N7531_2,
N7531_3,
N7531_4,
N7537_0,
N7537_1,
N7537_2,
N7537_3,
N7537_4,
N7543_0,
N7543_1,
N7543_2,
N7543_3,
N7543_4,
N7549_0,
N7549_1,
N7549_2,
N7549_3,
N7549_4,
N7555_0,
N7555_1,
N7555_2,
N7555_3,
N7555_4,
N7561_0,
N7561_1,
N7561_2,
N7561_3,
N7561_4,
N7567_0,
N7567_1,
N7567_2,
N7567_3,
N7567_4,
N7573_0,
N7573_1,
N7573_2,
N7573_3,
N7573_4,
N7579_0,
N7579_1,
N7582_0,
N7582_1,
N7589_0,
N7589_1,
N7592_0,
N7592_1,
N7595_0,
N7595_1,
N7712_0,
N7712_1,
N7715_0,
N7715_1,
N7724_0,
N7724_1,
N7762_0,
N7762_1,
N7765_0,
N7765_1,
N7772_0,
N7772_1,
N7775_0,
N7775_1,
N7778_0,
N7778_1,
N7800_0,
N7800_1,
N7803_0,
N7803_1,
N7812_0,
N7812_1,
N7826_0,
N7826_1,
N7829_0,
N7829_1,
N7836_0,
N7836_1,
N7839_0,
N7839_1,
N7842_0,
N7842_1,
N7864_0,
N7864_1,
N7867_0,
N7867_1,
N7876_0,
N7876_1,
N7890_0,
N7890_1,
N7893_0,
N7893_1,
N7900_0,
N7900_1,
N7903_0,
N7903_1,
N7906_0,
N7906_1,
N7932_0,
N7932_1,
N7935_0,
N7935_1,
N7940_0,
N7940_1,
N7954_0,
N7954_1,
N7957_0,
N7957_1,
N7960_0,
N7960_1,
N7963_0,
N7963_1,
N7970_0,
N7970_1,
N7998_0,
N7998_1,
N8001_0,
N8001_1,
N8004_0,
N8004_1,
N8013_0,
N8013_1,
N8017_0,
N8017_1,
N8045_0,
N8045_1,
N8048_0,
N8048_1,
N8061_0,
N8061_1,
N8064_0,
N8064_1,
N8079_0,
N8079_1,
N8082_0,
N8082_1,
N8093_0,
N8093_1,
N8096_0,
N8096_1,
N8099_0,
N8099_1,
N8102_0,
N8102_1;

fanout_n #(2, 0, 0) FANOUT_1 (N1, {N1_0, N1_1});
fanout_n #(6, 0, 0) FANOUT_2 (N4, {N4_0, N4_1, N4_2, N4_3, N4_4, N4_5});
fanout_n #(2, 0, 0) FANOUT_3 (N11, {N11_0, N11_1});
fanout_n #(2, 0, 0) FANOUT_4 (N14, {N14_0, N14_1});
fanout_n #(2, 0, 0) FANOUT_5 (N17, {N17_0, N17_1});
fanout_n #(2, 0, 0) FANOUT_6 (N20, {N20_0, N20_1});
fanout_n #(3, 0, 0) FANOUT_7 (N27, {N27_0, N27_1, N27_2});
fanout_n #(2, 0, 0) FANOUT_8 (N31, {N31_0, N31_1});
fanout_n #(2, 0, 0) FANOUT_9 (N34, {N34_0, N34_1});
fanout_n #(2, 0, 0) FANOUT_10 (N37, {N37_0, N37_1});
fanout_n #(2, 0, 0) FANOUT_11 (N40, {N40_0, N40_1});
fanout_n #(2, 0, 0) FANOUT_12 (N43, {N43_0, N43_1});
fanout_n #(2, 0, 0) FANOUT_13 (N46, {N46_0, N46_1});
fanout_n #(2, 0, 0) FANOUT_14 (N49, {N49_0, N49_1});
fanout_n #(6, 0, 0) FANOUT_15 (N54, {N54_0, N54_1, N54_2, N54_3, N54_4, N54_5});
fanout_n #(2, 0, 0) FANOUT_16 (N61, {N61_0, N61_1});
fanout_n #(2, 0, 0) FANOUT_17 (N64, {N64_0, N64_1});
fanout_n #(2, 0, 0) FANOUT_18 (N67, {N67_0, N67_1});
fanout_n #(2, 0, 0) FANOUT_19 (N70, {N70_0, N70_1});
fanout_n #(2, 0, 0) FANOUT_20 (N73, {N73_0, N73_1});
fanout_n #(2, 0, 0) FANOUT_21 (N76, {N76_0, N76_1});
fanout_n #(2, 0, 0) FANOUT_22 (N83, {N83_0, N83_1});
fanout_n #(2, 0, 0) FANOUT_23 (N88, {N88_0, N88_1});
fanout_n #(2, 0, 0) FANOUT_24 (N91, {N91_0, N91_1});
fanout_n #(2, 0, 0) FANOUT_25 (N94, {N94_0, N94_1});
fanout_n #(2, 0, 0) FANOUT_26 (N97, {N97_0, N97_1});
fanout_n #(2, 0, 0) FANOUT_27 (N100, {N100_0, N100_1});
fanout_n #(2, 0, 0) FANOUT_28 (N103, {N103_0, N103_1});
fanout_n #(2, 0, 0) FANOUT_29 (N106, {N106_0, N106_1});
fanout_n #(2, 0, 0) FANOUT_30 (N109, {N109_0, N109_1});
fanout_n #(2, 0, 0) FANOUT_31 (N123, {N123_0, N123_1});
fanout_n #(2, 0, 0) FANOUT_32 (N132, {N132_0, N132_1});
fanout_n #(2, 0, 0) FANOUT_33 (N137, {N137_0, N137_1});
fanout_n #(3, 0, 0) FANOUT_34 (N141, {N141_0, N141_1, N141_2});
fanout_n #(2, 0, 0) FANOUT_35 (N146, {N146_0, N146_1});
fanout_n #(2, 0, 0) FANOUT_36 (N149, {N149_0, N149_1});
fanout_n #(2, 0, 0) FANOUT_37 (N152, {N152_0, N152_1});
fanout_n #(2, 0, 0) FANOUT_38 (N155, {N155_0, N155_1});
fanout_n #(2, 0, 0) FANOUT_39 (N158, {N158_0, N158_1});
fanout_n #(2, 0, 0) FANOUT_40 (N161, {N161_0, N161_1});
fanout_n #(2, 0, 0) FANOUT_41 (N164, {N164_0, N164_1});
fanout_n #(2, 0, 0) FANOUT_42 (N167, {N167_0, N167_1});
fanout_n #(2, 0, 0) FANOUT_43 (N170, {N170_0, N170_1});
fanout_n #(2, 0, 0) FANOUT_44 (N173, {N173_0, N173_1});
fanout_n #(2, 0, 0) FANOUT_45 (N176, {N176_0, N176_1});
fanout_n #(2, 0, 0) FANOUT_46 (N179, {N179_0, N179_1});
fanout_n #(2, 0, 0) FANOUT_47 (N182, {N182_0, N182_1});
fanout_n #(2, 0, 0) FANOUT_48 (N185, {N185_0, N185_1});
fanout_n #(2, 0, 0) FANOUT_49 (N188, {N188_0, N188_1});
fanout_n #(2, 0, 0) FANOUT_50 (N191, {N191_0, N191_1});
fanout_n #(2, 0, 0) FANOUT_51 (N194, {N194_0, N194_1});
fanout_n #(2, 0, 0) FANOUT_52 (N197, {N197_0, N197_1});
fanout_n #(2, 0, 0) FANOUT_53 (N200, {N200_0, N200_1});
fanout_n #(2, 0, 0) FANOUT_54 (N203, {N203_0, N203_1});
fanout_n #(2, 0, 0) FANOUT_55 (N206, {N206_0, N206_1});
fanout_n #(6, 0, 0) FANOUT_56 (N210, {N210_0, N210_1, N210_2, N210_3, N210_4, N210_5});
fanout_n #(6, 0, 0) FANOUT_57 (N218, {N218_0, N218_1, N218_2, N218_3, N218_4, N218_5});
fanout_n #(6, 0, 0) FANOUT_58 (N226, {N226_0, N226_1, N226_2, N226_3, N226_4, N226_5});
fanout_n #(6, 0, 0) FANOUT_59 (N234, {N234_0, N234_1, N234_2, N234_3, N234_4, N234_5});
fanout_n #(2, 0, 0) FANOUT_60 (N242, {N242_0, N242_1});
fanout_n #(2, 0, 0) FANOUT_61 (N245, {N245_0, N245_1});
fanout_n #(2, 0, 0) FANOUT_62 (N248, {N248_0, N248_1});
fanout_n #(2, 0, 0) FANOUT_63 (N251, {N251_0, N251_1});
fanout_n #(2, 0, 0) FANOUT_64 (N254, {N254_0, N254_1});
fanout_n #(6, 0, 0) FANOUT_65 (N257, {N257_0, N257_1, N257_2, N257_3, N257_4, N257_5});
fanout_n #(6, 0, 0) FANOUT_66 (N265, {N265_0, N265_1, N265_2, N265_3, N265_4, N265_5});
fanout_n #(6, 0, 0) FANOUT_67 (N273, {N273_0, N273_1, N273_2, N273_3, N273_4, N273_5});
fanout_n #(6, 0, 0) FANOUT_68 (N281, {N281_0, N281_1, N281_2, N281_3, N281_4, N281_5});
fanout_n #(2, 0, 0) FANOUT_69 (N289, {N289_0, N289_1});
fanout_n #(5, 0, 0) FANOUT_70 (N293, {N293_0, N293_1, N293_2, N293_3, N293_4});
fanout_n #(2, 0, 0) FANOUT_71 (N299, {N299_0, N299_1});
fanout_n #(4, 0, 0) FANOUT_72 (N302, {N302_0, N302_1, N302_2, N302_3});
fanout_n #(6, 0, 0) FANOUT_73 (N308, {N308_0, N308_1, N308_2, N308_3, N308_4, N308_5});
fanout_n #(6, 0, 0) FANOUT_74 (N316, {N316_0, N316_1, N316_2, N316_3, N316_4, N316_5});
fanout_n #(6, 0, 0) FANOUT_75 (N324, {N324_0, N324_1, N324_2, N324_3, N324_4, N324_5});
fanout_n #(2, 0, 0) FANOUT_76 (N332, {N332_0, N332_1});
fanout_n #(2, 0, 0) FANOUT_77 (N335, {N335_0, N335_1});
fanout_n #(2, 0, 0) FANOUT_78 (N338, {N338_0, N338_1});
fanout_n #(6, 0, 0) FANOUT_79 (N341, {N341_0, N341_1, N341_2, N341_3, N341_4, N341_5});
fanout_n #(2, 0, 0) FANOUT_80 (N348, {N348_0, N348_1});
fanout_n #(6, 0, 0) FANOUT_81 (N351, {N351_0, N351_1, N351_2, N351_3, N351_4, N351_5});
fanout_n #(2, 0, 0) FANOUT_82 (N358, {N358_0, N358_1});
fanout_n #(4, 0, 0) FANOUT_83 (N361, {N361_0, N361_1, N361_2, N361_3});
fanout_n #(2, 0, 0) FANOUT_84 (N366, {N366_0, N366_1});
fanout_n #(2, 0, 0) FANOUT_85 (N369, {N369_0, N369_1});
fanout_n #(11, 0, 0) FANOUT_86 (N374, {N374_0, N374_1, N374_2, N374_3, N374_4, N374_5, N374_6, N374_7, N374_8, N374_9, N374_10});
fanout_n #(2, 0, 0) FANOUT_87 (N386, {N386_0, N386_1});
fanout_n #(10, 0, 0) FANOUT_88 (N389, {N389_0, N389_1, N389_2, N389_3, N389_4, N389_5, N389_6, N389_7, N389_8, N389_9});
fanout_n #(10, 0, 0) FANOUT_89 (N400, {N400_0, N400_1, N400_2, N400_3, N400_4, N400_5, N400_6, N400_7, N400_8, N400_9});
fanout_n #(10, 0, 0) FANOUT_90 (N411, {N411_0, N411_1, N411_2, N411_3, N411_4, N411_5, N411_6, N411_7, N411_8, N411_9});
fanout_n #(12, 0, 0) FANOUT_91 (N422, {N422_0, N422_1, N422_2, N422_3, N422_4, N422_5, N422_6, N422_7, N422_8, N422_9, N422_10, N422_11});
fanout_n #(10, 0, 0) FANOUT_92 (N435, {N435_0, N435_1, N435_2, N435_3, N435_4, N435_5, N435_6, N435_7, N435_8, N435_9});
fanout_n #(10, 0, 0) FANOUT_93 (N446, {N446_0, N446_1, N446_2, N446_3, N446_4, N446_5, N446_6, N446_7, N446_8, N446_9});
fanout_n #(10, 0, 0) FANOUT_94 (N457, {N457_0, N457_1, N457_2, N457_3, N457_4, N457_5, N457_6, N457_7, N457_8, N457_9});
fanout_n #(10, 0, 0) FANOUT_95 (N468, {N468_0, N468_1, N468_2, N468_3, N468_4, N468_5, N468_6, N468_7, N468_8, N468_9});
fanout_n #(10, 0, 0) FANOUT_96 (N479, {N479_0, N479_1, N479_2, N479_3, N479_4, N479_5, N479_6, N479_7, N479_8, N479_9});
fanout_n #(12, 0, 0) FANOUT_97 (N490, {N490_0, N490_1, N490_2, N490_3, N490_4, N490_5, N490_6, N490_7, N490_8, N490_9, N490_10, N490_11});
fanout_n #(10, 0, 0) FANOUT_98 (N503, {N503_0, N503_1, N503_2, N503_3, N503_4, N503_5, N503_6, N503_7, N503_8, N503_9});
fanout_n #(8, 0, 0) FANOUT_99 (N514, {N514_0, N514_1, N514_2, N514_3, N514_4, N514_5, N514_6, N514_7});
fanout_n #(10, 0, 0) FANOUT_100 (N523, {N523_0, N523_1, N523_2, N523_3, N523_4, N523_5, N523_6, N523_7, N523_8, N523_9});
fanout_n #(10, 0, 0) FANOUT_101 (N534, {N534_0, N534_1, N534_2, N534_3, N534_4, N534_5, N534_6, N534_7, N534_8, N534_9});
fanout_n #(3, 0, 0) FANOUT_102 (N545, {N545_0, N545_1, N545_2});
fanout_n #(2, 0, 0) FANOUT_103 (N549, {N549_0, N549_1});
fanout_n #(3, 0, 0) FANOUT_104 (N552, {N552_0, N552_1, N552_2});
fanout_n #(2, 0, 0) FANOUT_105 (N556, {N556_0, N556_1});
fanout_n #(2, 0, 0) FANOUT_106 (N559, {N559_0, N559_1});
fanout_n #(3, 0, 0) FANOUT_107 (N562, {N562_0, N562_1, N562_2});
fanout_n #(4, 0, 0) FANOUT_108 (N566, {N566_0, N566_1, N566_2, N566_3});
fanout_n #(2, 0, 0) FANOUT_109 (N571, {N571_0, N571_1});
fanout_n #(2, 0, 0) FANOUT_110 (N574, {N574_0, N574_1});
fanout_n #(2, 0, 0) FANOUT_111 (N577, {N577_0, N577_1});
fanout_n #(2, 0, 0) FANOUT_112 (N580, {N580_0, N580_1});
fanout_n #(4, 0, 0) FANOUT_113 (N583, {N583_0, N583_1, N583_2, N583_3});
fanout_n #(2, 0, 0) FANOUT_114 (N588, {N588_0, N588_1});
fanout_n #(2, 0, 0) FANOUT_115 (N592, {N592_0, N592_1});
fanout_n #(3, 0, 0) FANOUT_116 (N599, {N599_0, N599_1, N599_2});
fanout_n #(3, 0, 0) FANOUT_117 (N603, {N603_0, N603_1, N603_2});
fanout_n #(2, 0, 0) FANOUT_118 (N607, {N607_0, N607_1});
fanout_n #(2, 0, 0) FANOUT_119 (N610, {N610_0, N610_1});
fanout_n #(2, 0, 0) FANOUT_120 (N613, {N613_0, N613_1});
fanout_n #(2, 0, 0) FANOUT_121 (N616, {N616_0, N616_1});
fanout_n #(5, 0, 0) FANOUT_122 (N619, {N619_0, N619_1, N619_2, N619_3, N619_4});
fanout_n #(5, 0, 0) FANOUT_123 (N625, {N625_0, N625_1, N625_2, N625_3, N625_4});
fanout_n #(12, 0, 0) FANOUT_124 (N1067, {N1067_0, N1067_1, N1067_2, N1067_3, N1067_4, N1067_5, N1067_6, N1067_7, N1067_8, N1067_9, N1067_10, N1067_11});
fanout_n #(11, 0, 0) FANOUT_125 (N1080, {N1080_0, N1080_1, N1080_2, N1080_3, N1080_4, N1080_5, N1080_6, N1080_7, N1080_8, N1080_9, N1080_10});
fanout_n #(11, 0, 0) FANOUT_126 (N1092, {N1092_0, N1092_1, N1092_2, N1092_3, N1092_4, N1092_5, N1092_6, N1092_7, N1092_8, N1092_9, N1092_10});
fanout_n #(12, 0, 0) FANOUT_127 (N1104, {N1104_0, N1104_1, N1104_2, N1104_3, N1104_4, N1104_5, N1104_6, N1104_7, N1104_8, N1104_9, N1104_10, N1104_11});
fanout_n #(3, 0, 0) FANOUT_128 (N1157, {N1157_0, N1157_1, N1157_2});
fanout_n #(11, 0, 0) FANOUT_129 (N1161, {N1161_0, N1161_1, N1161_2, N1161_3, N1161_4, N1161_5, N1161_6, N1161_7, N1161_8, N1161_9, N1161_10});
fanout_n #(11, 0, 0) FANOUT_130 (N1173, {N1173_0, N1173_1, N1173_2, N1173_3, N1173_4, N1173_5, N1173_6, N1173_7, N1173_8, N1173_9, N1173_10});
fanout_n #(11, 0, 0) FANOUT_131 (N1185, {N1185_0, N1185_1, N1185_2, N1185_3, N1185_4, N1185_5, N1185_6, N1185_7, N1185_8, N1185_9, N1185_10});
fanout_n #(11, 0, 0) FANOUT_132 (N1197, {N1197_0, N1197_1, N1197_2, N1197_3, N1197_4, N1197_5, N1197_6, N1197_7, N1197_8, N1197_9, N1197_10});
fanout_n #(3, 0, 0) FANOUT_133 (N1209, {N1209_0, N1209_1, N1209_2});
fanout_n #(2, 0, 0) FANOUT_134 (N1213, {N1213_0, N1213_1});
fanout_n #(2, 0, 0) FANOUT_135 (N1216, {N1216_0, N1216_1});
fanout_n #(3, 0, 0) FANOUT_136 (N1219, {N1219_0, N1219_1, N1219_2});
fanout_n #(11, 0, 0) FANOUT_137 (N1223, {N1223_0, N1223_1, N1223_2, N1223_3, N1223_4, N1223_5, N1223_6, N1223_7, N1223_8, N1223_9, N1223_10});
fanout_n #(11, 0, 0) FANOUT_138 (N1235, {N1235_0, N1235_1, N1235_2, N1235_3, N1235_4, N1235_5, N1235_6, N1235_7, N1235_8, N1235_9, N1235_10});
fanout_n #(11, 0, 0) FANOUT_139 (N1247, {N1247_0, N1247_1, N1247_2, N1247_3, N1247_4, N1247_5, N1247_6, N1247_7, N1247_8, N1247_9, N1247_10});
fanout_n #(11, 0, 0) FANOUT_140 (N1259, {N1259_0, N1259_1, N1259_2, N1259_3, N1259_4, N1259_5, N1259_6, N1259_7, N1259_8, N1259_9, N1259_10});
fanout_n #(8, 0, 0) FANOUT_141 (N1271, {N1271_0, N1271_1, N1271_2, N1271_3, N1271_4, N1271_5, N1271_6, N1271_7});
fanout_n #(11, 0, 0) FANOUT_142 (N1280, {N1280_0, N1280_1, N1280_2, N1280_3, N1280_4, N1280_5, N1280_6, N1280_7, N1280_8, N1280_9, N1280_10});
fanout_n #(10, 0, 0) FANOUT_143 (N1292, {N1292_0, N1292_1, N1292_2, N1292_3, N1292_4, N1292_5, N1292_6, N1292_7, N1292_8, N1292_9});
fanout_n #(11, 0, 0) FANOUT_144 (N1303, {N1303_0, N1303_1, N1303_2, N1303_3, N1303_4, N1303_5, N1303_6, N1303_7, N1303_8, N1303_9, N1303_10});
fanout_n #(11, 0, 0) FANOUT_145 (N1315, {N1315_0, N1315_1, N1315_2, N1315_3, N1315_4, N1315_5, N1315_6, N1315_7, N1315_8, N1315_9, N1315_10});
fanout_n #(11, 0, 0) FANOUT_146 (N1327, {N1327_0, N1327_1, N1327_2, N1327_3, N1327_4, N1327_5, N1327_6, N1327_7, N1327_8, N1327_9, N1327_10});
fanout_n #(11, 0, 0) FANOUT_147 (N1339, {N1339_0, N1339_1, N1339_2, N1339_3, N1339_4, N1339_5, N1339_6, N1339_7, N1339_8, N1339_9, N1339_10});
fanout_n #(11, 0, 0) FANOUT_148 (N1351, {N1351_0, N1351_1, N1351_2, N1351_3, N1351_4, N1351_5, N1351_6, N1351_7, N1351_8, N1351_9, N1351_10});
fanout_n #(11, 0, 0) FANOUT_149 (N1363, {N1363_0, N1363_1, N1363_2, N1363_3, N1363_4, N1363_5, N1363_6, N1363_7, N1363_8, N1363_9, N1363_10});
fanout_n #(2, 0, 0) FANOUT_150 (N1375, {N1375_0, N1375_1});
fanout_n #(2, 0, 0) FANOUT_151 (N1378, {N1378_0, N1378_1});
fanout_n #(2, 0, 0) FANOUT_152 (N1381, {N1381_0, N1381_1});
fanout_n #(2, 0, 0) FANOUT_153 (N1384, {N1384_0, N1384_1});
fanout_n #(2, 0, 0) FANOUT_154 (N1387, {N1387_0, N1387_1});
fanout_n #(2, 0, 0) FANOUT_155 (N1390, {N1390_0, N1390_1});
fanout_n #(2, 0, 0) FANOUT_156 (N1393, {N1393_0, N1393_1});
fanout_n #(2, 0, 0) FANOUT_157 (N1396, {N1396_0, N1396_1});
fanout_n #(2, 0, 0) FANOUT_158 (N1415, {N1415_0, N1415_1});
fanout_n #(2, 0, 0) FANOUT_159 (N1418, {N1418_0, N1418_1});
fanout_n #(2, 0, 0) FANOUT_160 (N1421, {N1421_0, N1421_1});
fanout_n #(2, 0, 0) FANOUT_161 (N1424, {N1424_0, N1424_1});
fanout_n #(2, 0, 0) FANOUT_162 (N1427, {N1427_0, N1427_1});
fanout_n #(2, 0, 0) FANOUT_163 (N1430, {N1430_0, N1430_1});
fanout_n #(2, 0, 0) FANOUT_164 (N1433, {N1433_0, N1433_1});
fanout_n #(2, 0, 0) FANOUT_165 (N1436, {N1436_0, N1436_1});
fanout_n #(6, 0, 0) FANOUT_166 (N1455, {N1455_0, N1455_1, N1455_2, N1455_3, N1455_4, N1455_5});
fanout_n #(6, 0, 0) FANOUT_167 (N1462, {N1462_0, N1462_1, N1462_2, N1462_3, N1462_4, N1462_5});
fanout_n #(5, 0, 0) FANOUT_168 (N1469, {N1469_0, N1469_1, N1469_2, N1469_3, N1469_4});
fanout_n #(3, 0, 0) FANOUT_169 (N1475, {N1475_0, N1475_1, N1475_2});
fanout_n #(2, 0, 0) FANOUT_170 (N1479, {N1479_0, N1479_1});
fanout_n #(9, 0, 0) FANOUT_171 (N1482, {N1482_0, N1482_1, N1482_2, N1482_3, N1482_4, N1482_5, N1482_6, N1482_7, N1482_8});
fanout_n #(2, 0, 0) FANOUT_172 (N1492, {N1492_0, N1492_1});
fanout_n #(2, 0, 0) FANOUT_173 (N1495, {N1495_0, N1495_1});
fanout_n #(2, 0, 0) FANOUT_174 (N1498, {N1498_0, N1498_1});
fanout_n #(2, 0, 0) FANOUT_175 (N1501, {N1501_0, N1501_1});
fanout_n #(2, 0, 0) FANOUT_176 (N1504, {N1504_0, N1504_1});
fanout_n #(2, 0, 0) FANOUT_177 (N1507, {N1507_0, N1507_1});
fanout_n #(2, 0, 0) FANOUT_178 (N1510, {N1510_0, N1510_1});
fanout_n #(2, 0, 0) FANOUT_179 (N1513, {N1513_0, N1513_1});
fanout_n #(2, 0, 0) FANOUT_180 (N1516, {N1516_0, N1516_1});
fanout_n #(2, 0, 0) FANOUT_181 (N1519, {N1519_0, N1519_1});
fanout_n #(2, 0, 0) FANOUT_182 (N1522, {N1522_0, N1522_1});
fanout_n #(2, 0, 0) FANOUT_183 (N1525, {N1525_0, N1525_1});
fanout_n #(2, 0, 0) FANOUT_184 (N1542, {N1542_0, N1542_1});
fanout_n #(2, 0, 0) FANOUT_185 (N1545, {N1545_0, N1545_1});
fanout_n #(2, 0, 0) FANOUT_186 (N1548, {N1548_0, N1548_1});
fanout_n #(2, 0, 0) FANOUT_187 (N1551, {N1551_0, N1551_1});
fanout_n #(2, 0, 0) FANOUT_188 (N1554, {N1554_0, N1554_1});
fanout_n #(2, 0, 0) FANOUT_189 (N1557, {N1557_0, N1557_1});
fanout_n #(2, 0, 0) FANOUT_190 (N1560, {N1560_0, N1560_1});
fanout_n #(2, 0, 0) FANOUT_191 (N1563, {N1563_0, N1563_1});
fanout_n #(6, 0, 0) FANOUT_192 (N1566, {N1566_0, N1566_1, N1566_2, N1566_3, N1566_4, N1566_5});
fanout_n #(6, 0, 0) FANOUT_193 (N1573, {N1573_0, N1573_1, N1573_2, N1573_3, N1573_4, N1573_5});
fanout_n #(2, 0, 0) FANOUT_194 (N1580, {N1580_0, N1580_1});
fanout_n #(4, 0, 0) FANOUT_195 (N1583, {N1583_0, N1583_1, N1583_2, N1583_3});
fanout_n #(5, 0, 0) FANOUT_196 (N1588, {N1588_0, N1588_1, N1588_2, N1588_3, N1588_4});
fanout_n #(2, 0, 0) FANOUT_197 (N1594, {N1594_0, N1594_1});
fanout_n #(2, 0, 0) FANOUT_198 (N1597, {N1597_0, N1597_1});
fanout_n #(2, 0, 0) FANOUT_199 (N1600, {N1600_0, N1600_1});
fanout_n #(2, 0, 0) FANOUT_200 (N1603, {N1603_0, N1603_1});
fanout_n #(2, 0, 0) FANOUT_201 (N1606, {N1606_0, N1606_1});
fanout_n #(2, 0, 0) FANOUT_202 (N1609, {N1609_0, N1609_1});
fanout_n #(2, 0, 0) FANOUT_203 (N1612, {N1612_0, N1612_1});
fanout_n #(2, 0, 0) FANOUT_204 (N1615, {N1615_0, N1615_1});
fanout_n #(2, 0, 0) FANOUT_205 (N1618, {N1618_0, N1618_1});
fanout_n #(2, 0, 0) FANOUT_206 (N1621, {N1621_0, N1621_1});
fanout_n #(2, 0, 0) FANOUT_207 (N1624, {N1624_0, N1624_1});
fanout_n #(2, 0, 0) FANOUT_208 (N1627, {N1627_0, N1627_1});
fanout_n #(2, 0, 0) FANOUT_209 (N1630, {N1630_0, N1630_1});
fanout_n #(2, 0, 0) FANOUT_210 (N1633, {N1633_0, N1633_1});
fanout_n #(2, 0, 0) FANOUT_211 (N1636, {N1636_0, N1636_1});
fanout_n #(2, 0, 0) FANOUT_212 (N1639, {N1639_0, N1639_1});
fanout_n #(2, 0, 0) FANOUT_213 (N1642, {N1642_0, N1642_1});
fanout_n #(2, 0, 0) FANOUT_214 (N1645, {N1645_0, N1645_1});
fanout_n #(2, 0, 0) FANOUT_215 (N1648, {N1648_0, N1648_1});
fanout_n #(2, 0, 0) FANOUT_216 (N1651, {N1651_0, N1651_1});
fanout_n #(2, 0, 0) FANOUT_217 (N1654, {N1654_0, N1654_1});
fanout_n #(2, 0, 0) FANOUT_218 (N1657, {N1657_0, N1657_1});
fanout_n #(2, 0, 0) FANOUT_219 (N1660, {N1660_0, N1660_1});
fanout_n #(11, 0, 0) FANOUT_220 (N1663, {N1663_0, N1663_1, N1663_2, N1663_3, N1663_4, N1663_5, N1663_6, N1663_7, N1663_8, N1663_9, N1663_10});
fanout_n #(9, 0, 0) FANOUT_221 (N1675, {N1675_0, N1675_1, N1675_2, N1675_3, N1675_4, N1675_5, N1675_6, N1675_7, N1675_8});
fanout_n #(11, 0, 0) FANOUT_222 (N1685, {N1685_0, N1685_1, N1685_2, N1685_3, N1685_4, N1685_5, N1685_6, N1685_7, N1685_8, N1685_9, N1685_10});
fanout_n #(11, 0, 0) FANOUT_223 (N1697, {N1697_0, N1697_1, N1697_2, N1697_3, N1697_4, N1697_5, N1697_6, N1697_7, N1697_8, N1697_9, N1697_10});
fanout_n #(11, 0, 0) FANOUT_224 (N1709, {N1709_0, N1709_1, N1709_2, N1709_3, N1709_4, N1709_5, N1709_6, N1709_7, N1709_8, N1709_9, N1709_10});
fanout_n #(5, 0, 0) FANOUT_225 (N1721, {N1721_0, N1721_1, N1721_2, N1721_3, N1721_4});
fanout_n #(3, 0, 0) FANOUT_226 (N1727, {N1727_0, N1727_1, N1727_2});
fanout_n #(11, 0, 0) FANOUT_227 (N1731, {N1731_0, N1731_1, N1731_2, N1731_3, N1731_4, N1731_5, N1731_6, N1731_7, N1731_8, N1731_9, N1731_10});
fanout_n #(11, 0, 0) FANOUT_228 (N1743, {N1743_0, N1743_1, N1743_2, N1743_3, N1743_4, N1743_5, N1743_6, N1743_7, N1743_8, N1743_9, N1743_10});
fanout_n #(2, 0, 0) FANOUT_229 (N1755, {N1755_0, N1755_1});
fanout_n #(2, 0, 0) FANOUT_230 (N1758, {N1758_0, N1758_1});
fanout_n #(7, 0, 0) FANOUT_231 (N1761, {N1761_0, N1761_1, N1761_2, N1761_3, N1761_4, N1761_5, N1761_6});
fanout_n #(7, 0, 0) FANOUT_232 (N1769, {N1769_0, N1769_1, N1769_2, N1769_3, N1769_4, N1769_5, N1769_6});
fanout_n #(7, 0, 0) FANOUT_233 (N1777, {N1777_0, N1777_1, N1777_2, N1777_3, N1777_4, N1777_5, N1777_6});
fanout_n #(7, 0, 0) FANOUT_234 (N1785, {N1785_0, N1785_1, N1785_2, N1785_3, N1785_4, N1785_5, N1785_6});
fanout_n #(6, 0, 0) FANOUT_235 (N1793, {N1793_0, N1793_1, N1793_2, N1793_3, N1793_4, N1793_5});
fanout_n #(6, 0, 0) FANOUT_236 (N1800, {N1800_0, N1800_1, N1800_2, N1800_3, N1800_4, N1800_5});
fanout_n #(6, 0, 0) FANOUT_237 (N1807, {N1807_0, N1807_1, N1807_2, N1807_3, N1807_4, N1807_5});
fanout_n #(6, 0, 0) FANOUT_238 (N1814, {N1814_0, N1814_1, N1814_2, N1814_3, N1814_4, N1814_5});
fanout_n #(2, 0, 0) FANOUT_239 (N1821, {N1821_0, N1821_1});
fanout_n #(2, 0, 0) FANOUT_240 (N1824, {N1824_0, N1824_1});
fanout_n #(2, 0, 0) FANOUT_241 (N1827, {N1827_0, N1827_1});
fanout_n #(2, 0, 0) FANOUT_242 (N1830, {N1830_0, N1830_1});
fanout_n #(2, 0, 0) FANOUT_243 (N1833, {N1833_0, N1833_1});
fanout_n #(2, 0, 0) FANOUT_244 (N1836, {N1836_0, N1836_1});
fanout_n #(2, 0, 0) FANOUT_245 (N1839, {N1839_0, N1839_1});
fanout_n #(2, 0, 0) FANOUT_246 (N1842, {N1842_0, N1842_1});
fanout_n #(2, 0, 0) FANOUT_247 (N1845, {N1845_0, N1845_1});
fanout_n #(2, 0, 0) FANOUT_248 (N1848, {N1848_0, N1848_1});
fanout_n #(2, 0, 0) FANOUT_249 (N1851, {N1851_0, N1851_1});
fanout_n #(2, 0, 0) FANOUT_250 (N1854, {N1854_0, N1854_1});
fanout_n #(2, 0, 0) FANOUT_251 (N1857, {N1857_0, N1857_1});
fanout_n #(2, 0, 0) FANOUT_252 (N1860, {N1860_0, N1860_1});
fanout_n #(2, 0, 0) FANOUT_253 (N1863, {N1863_0, N1863_1});
fanout_n #(2, 0, 0) FANOUT_254 (N1866, {N1866_0, N1866_1});
fanout_n #(2, 0, 0) FANOUT_255 (N1869, {N1869_0, N1869_1});
fanout_n #(2, 0, 0) FANOUT_256 (N1872, {N1872_0, N1872_1});
fanout_n #(2, 0, 0) FANOUT_257 (N1875, {N1875_0, N1875_1});
fanout_n #(2, 0, 0) FANOUT_258 (N1878, {N1878_0, N1878_1});
fanout_n #(2, 0, 0) FANOUT_259 (N1881, {N1881_0, N1881_1});
fanout_n #(2, 0, 0) FANOUT_260 (N1884, {N1884_0, N1884_1});
fanout_n #(2, 0, 0) FANOUT_261 (N1887, {N1887_0, N1887_1});
fanout_n #(2, 0, 0) FANOUT_262 (N1890, {N1890_0, N1890_1});
fanout_n #(2, 0, 0) FANOUT_263 (N1893, {N1893_0, N1893_1});
fanout_n #(2, 0, 0) FANOUT_264 (N1896, {N1896_0, N1896_1});
fanout_n #(2, 0, 0) FANOUT_265 (N1899, {N1899_0, N1899_1});
fanout_n #(2, 0, 0) FANOUT_266 (N1902, {N1902_0, N1902_1});
fanout_n #(2, 0, 0) FANOUT_267 (N1905, {N1905_0, N1905_1});
fanout_n #(2, 0, 0) FANOUT_268 (N1908, {N1908_0, N1908_1});
fanout_n #(2, 0, 0) FANOUT_269 (N1911, {N1911_0, N1911_1});
fanout_n #(2, 0, 0) FANOUT_270 (N1914, {N1914_0, N1914_1});
fanout_n #(2, 0, 0) FANOUT_271 (N1917, {N1917_0, N1917_1});
fanout_n #(2, 0, 0) FANOUT_272 (N1920, {N1920_0, N1920_1});
fanout_n #(2, 0, 0) FANOUT_273 (N1923, {N1923_0, N1923_1});
fanout_n #(2, 0, 0) FANOUT_274 (N1926, {N1926_0, N1926_1});
fanout_n #(2, 0, 0) FANOUT_275 (N1929, {N1929_0, N1929_1});
fanout_n #(2, 0, 0) FANOUT_276 (N1932, {N1932_0, N1932_1});
fanout_n #(2, 0, 0) FANOUT_277 (N1935, {N1935_0, N1935_1});
fanout_n #(2, 0, 0) FANOUT_278 (N1938, {N1938_0, N1938_1});
fanout_n #(2, 0, 0) FANOUT_279 (N1941, {N1941_0, N1941_1});
fanout_n #(2, 0, 0) FANOUT_280 (N1944, {N1944_0, N1944_1});
fanout_n #(2, 0, 0) FANOUT_281 (N1947, {N1947_0, N1947_1});
fanout_n #(2, 0, 0) FANOUT_282 (N1950, {N1950_0, N1950_1});
fanout_n #(2, 0, 0) FANOUT_283 (N1953, {N1953_0, N1953_1});
fanout_n #(2, 0, 0) FANOUT_284 (N1956, {N1956_0, N1956_1});
fanout_n #(2, 0, 0) FANOUT_285 (N1959, {N1959_0, N1959_1});
fanout_n #(2, 0, 0) FANOUT_286 (N1962, {N1962_0, N1962_1});
fanout_n #(2, 0, 0) FANOUT_287 (N1965, {N1965_0, N1965_1});
fanout_n #(2, 0, 0) FANOUT_288 (N1968, {N1968_0, N1968_1});
fanout_n #(5, 0, 0) FANOUT_289 (N2647, {N2647_0, N2647_1, N2647_2, N2647_3, N2647_4});
fanout_n #(10, 0, 0) FANOUT_290 (N2653, {N2653_0, N2653_1, N2653_2, N2653_3, N2653_4, N2653_5, N2653_6, N2653_7, N2653_8, N2653_9});
fanout_n #(10, 0, 0) FANOUT_291 (N2664, {N2664_0, N2664_1, N2664_2, N2664_3, N2664_4, N2664_5, N2664_6, N2664_7, N2664_8, N2664_9});
fanout_n #(5, 0, 0) FANOUT_292 (N2675, {N2675_0, N2675_1, N2675_2, N2675_3, N2675_4});
fanout_n #(10, 0, 0) FANOUT_293 (N2681, {N2681_0, N2681_1, N2681_2, N2681_3, N2681_4, N2681_5, N2681_6, N2681_7, N2681_8, N2681_9});
fanout_n #(10, 0, 0) FANOUT_294 (N2692, {N2692_0, N2692_1, N2692_2, N2692_3, N2692_4, N2692_5, N2692_6, N2692_7, N2692_8, N2692_9});
fanout_n #(4, 0, 0) FANOUT_295 (N2704, {N2704_0, N2704_1, N2704_2, N2704_3});
fanout_n #(5, 0, 0) FANOUT_296 (N2722, {N2722_0, N2722_1, N2722_2, N2722_3, N2722_4});
fanout_n #(10, 0, 0) FANOUT_297 (N2728, {N2728_0, N2728_1, N2728_2, N2728_3, N2728_4, N2728_5, N2728_6, N2728_7, N2728_8, N2728_9});
fanout_n #(10, 0, 0) FANOUT_298 (N2739, {N2739_0, N2739_1, N2739_2, N2739_3, N2739_4, N2739_5, N2739_6, N2739_7, N2739_8, N2739_9});
fanout_n #(5, 0, 0) FANOUT_299 (N2750, {N2750_0, N2750_1, N2750_2, N2750_3, N2750_4});
fanout_n #(10, 0, 0) FANOUT_300 (N2756, {N2756_0, N2756_1, N2756_2, N2756_3, N2756_4, N2756_5, N2756_6, N2756_7, N2756_8, N2756_9});
fanout_n #(10, 0, 0) FANOUT_301 (N2767, {N2767_0, N2767_1, N2767_2, N2767_3, N2767_4, N2767_5, N2767_6, N2767_7, N2767_8, N2767_9});
fanout_n #(10, 0, 0) FANOUT_302 (N2779, {N2779_0, N2779_1, N2779_2, N2779_3, N2779_4, N2779_5, N2779_6, N2779_7, N2779_8, N2779_9});
fanout_n #(10, 0, 0) FANOUT_303 (N2790, {N2790_0, N2790_1, N2790_2, N2790_3, N2790_4, N2790_5, N2790_6, N2790_7, N2790_8, N2790_9});
fanout_n #(10, 0, 0) FANOUT_304 (N2801, {N2801_0, N2801_1, N2801_2, N2801_3, N2801_4, N2801_5, N2801_6, N2801_7, N2801_8, N2801_9});
fanout_n #(10, 0, 0) FANOUT_305 (N2812, {N2812_0, N2812_1, N2812_2, N2812_3, N2812_4, N2812_5, N2812_6, N2812_7, N2812_8, N2812_9});
fanout_n #(5, 0, 0) FANOUT_306 (N2855, {N2855_0, N2855_1, N2855_2, N2855_3, N2855_4});
fanout_n #(5, 0, 0) FANOUT_307 (N2861, {N2861_0, N2861_1, N2861_2, N2861_3, N2861_4});
fanout_n #(4, 0, 0) FANOUT_308 (N2877, {N2877_0, N2877_1, N2877_2, N2877_3});
fanout_n #(8, 0, 0) FANOUT_309 (N2882, {N2882_0, N2882_1, N2882_2, N2882_3, N2882_4, N2882_5, N2882_6, N2882_7});
fanout_n #(9, 0, 0) FANOUT_310 (N2891, {N2891_0, N2891_1, N2891_2, N2891_3, N2891_4, N2891_5, N2891_6, N2891_7, N2891_8});
fanout_n #(5, 0, 0) FANOUT_311 (N2942, {N2942_0, N2942_1, N2942_2, N2942_3, N2942_4});
fanout_n #(5, 0, 0) FANOUT_312 (N2948, {N2948_0, N2948_1, N2948_2, N2948_3, N2948_4});
fanout_n #(4, 0, 0) FANOUT_313 (N2964, {N2964_0, N2964_1, N2964_2, N2964_3});
fanout_n #(2, 0, 0) FANOUT_314 (N3000, {N3000_0, N3000_1});
fanout_n #(2, 0, 0) FANOUT_315 (N3003, {N3003_0, N3003_1});
fanout_n #(2, 0, 0) FANOUT_316 (N3007, {N3007_0, N3007_1});
fanout_n #(2, 0, 0) FANOUT_317 (N3010, {N3010_0, N3010_1});
fanout_n #(2, 0, 0) FANOUT_318 (N3035, {N3035_0, N3035_1});
fanout_n #(2, 0, 0) FANOUT_319 (N3038, {N3038_0, N3038_1});
fanout_n #(10, 0, 0) FANOUT_320 (N3041, {N3041_0, N3041_1, N3041_2, N3041_3, N3041_4, N3041_5, N3041_6, N3041_7, N3041_8, N3041_9});
fanout_n #(10, 0, 0) FANOUT_321 (N3052, {N3052_0, N3052_1, N3052_2, N3052_3, N3052_4, N3052_5, N3052_6, N3052_7, N3052_8, N3052_9});
fanout_n #(4, 0, 0) FANOUT_322 (N3063, {N3063_0, N3063_1, N3063_2, N3063_3});
fanout_n #(2, 0, 0) FANOUT_323 (N3068, {N3068_0, N3068_1});
fanout_n #(10, 0, 0) FANOUT_324 (N3075, {N3075_0, N3075_1, N3075_2, N3075_3, N3075_4, N3075_5, N3075_6, N3075_7, N3075_8, N3075_9});
fanout_n #(10, 0, 0) FANOUT_325 (N3086, {N3086_0, N3086_1, N3086_2, N3086_3, N3086_4, N3086_5, N3086_6, N3086_7, N3086_8, N3086_9});
fanout_n #(10, 0, 0) FANOUT_326 (N3097, {N3097_0, N3097_1, N3097_2, N3097_3, N3097_4, N3097_5, N3097_6, N3097_7, N3097_8, N3097_9});
fanout_n #(10, 0, 0) FANOUT_327 (N3108, {N3108_0, N3108_1, N3108_2, N3108_3, N3108_4, N3108_5, N3108_6, N3108_7, N3108_8, N3108_9});
fanout_n #(10, 0, 0) FANOUT_328 (N3119, {N3119_0, N3119_1, N3119_2, N3119_3, N3119_4, N3119_5, N3119_6, N3119_7, N3119_8, N3119_9});
fanout_n #(10, 0, 0) FANOUT_329 (N3130, {N3130_0, N3130_1, N3130_2, N3130_3, N3130_4, N3130_5, N3130_6, N3130_7, N3130_8, N3130_9});
fanout_n #(10, 0, 0) FANOUT_330 (N3147, {N3147_0, N3147_1, N3147_2, N3147_3, N3147_4, N3147_5, N3147_6, N3147_7, N3147_8, N3147_9});
fanout_n #(10, 0, 0) FANOUT_331 (N3158, {N3158_0, N3158_1, N3158_2, N3158_3, N3158_4, N3158_5, N3158_6, N3158_7, N3158_8, N3158_9});
fanout_n #(10, 0, 0) FANOUT_332 (N3169, {N3169_0, N3169_1, N3169_2, N3169_3, N3169_4, N3169_5, N3169_6, N3169_7, N3169_8, N3169_9});
fanout_n #(10, 0, 0) FANOUT_333 (N3180, {N3180_0, N3180_1, N3180_2, N3180_3, N3180_4, N3180_5, N3180_6, N3180_7, N3180_8, N3180_9});
fanout_n #(2, 0, 0) FANOUT_334 (N3191, {N3191_0, N3191_1});
fanout_n #(2, 0, 0) FANOUT_335 (N3200, {N3200_0, N3200_1});
fanout_n #(2, 0, 0) FANOUT_336 (N3456, {N3456_0, N3456_1});
fanout_n #(8, 0, 0) FANOUT_337 (N3691, {N3691_0, N3691_1, N3691_2, N3691_3, N3691_4, N3691_5, N3691_6, N3691_7});
fanout_n #(2, 0, 0) FANOUT_338 (N3705, {N3705_0, N3705_1});
fanout_n #(5, 0, 0) FANOUT_339 (N3732, {N3732_0, N3732_1, N3732_2, N3732_3, N3732_4});
fanout_n #(3, 0, 0) FANOUT_340 (N3771, {N3771_0, N3771_1, N3771_2});
fanout_n #(3, 0, 0) FANOUT_341 (N3775, {N3775_0, N3775_1, N3775_2});
fanout_n #(3, 0, 0) FANOUT_342 (N3789, {N3789_0, N3789_1, N3789_2});
fanout_n #(3, 0, 0) FANOUT_343 (N3793, {N3793_0, N3793_1, N3793_2});
fanout_n #(2, 0, 0) FANOUT_344 (N3797, {N3797_0, N3797_1});
fanout_n #(2, 0, 0) FANOUT_345 (N3810, {N3810_0, N3810_1});
fanout_n #(2, 0, 0) FANOUT_346 (N3813, {N3813_0, N3813_1});
fanout_n #(2, 0, 0) FANOUT_347 (N3816, {N3816_0, N3816_1});
fanout_n #(2, 0, 0) FANOUT_348 (N3819, {N3819_0, N3819_1});
fanout_n #(2, 0, 0) FANOUT_349 (N3824, {N3824_0, N3824_1});
fanout_n #(6, 0, 0) FANOUT_350 (N3842, {N3842_0, N3842_1, N3842_2, N3842_3, N3842_4, N3842_5});
fanout_n #(5, 0, 0) FANOUT_351 (N3849, {N3849_0, N3849_1, N3849_2, N3849_3, N3849_4});
fanout_n #(5, 0, 0) FANOUT_352 (N3855, {N3855_0, N3855_1, N3855_2, N3855_3, N3855_4});
fanout_n #(5, 0, 0) FANOUT_353 (N3861, {N3861_0, N3861_1, N3861_2, N3861_3, N3861_4});
fanout_n #(5, 0, 0) FANOUT_354 (N3867, {N3867_0, N3867_1, N3867_2, N3867_3, N3867_4});
fanout_n #(7, 0, 0) FANOUT_355 (N3873, {N3873_0, N3873_1, N3873_2, N3873_3, N3873_4, N3873_5, N3873_6});
fanout_n #(5, 0, 0) FANOUT_356 (N3881, {N3881_0, N3881_1, N3881_2, N3881_3, N3881_4});
fanout_n #(5, 0, 0) FANOUT_357 (N3887, {N3887_0, N3887_1, N3887_2, N3887_3, N3887_4});
fanout_n #(5, 0, 0) FANOUT_358 (N3893, {N3893_0, N3893_1, N3893_2, N3893_3, N3893_4});
fanout_n #(2, 0, 0) FANOUT_359 (N3911, {N3911_0, N3911_1});
fanout_n #(5, 0, 0) FANOUT_360 (N3921, {N3921_0, N3921_1, N3921_2, N3921_3, N3921_4});
fanout_n #(5, 0, 0) FANOUT_361 (N3927, {N3927_0, N3927_1, N3927_2, N3927_3, N3927_4});
fanout_n #(5, 0, 0) FANOUT_362 (N3933, {N3933_0, N3933_1, N3933_2, N3933_3, N3933_4});
fanout_n #(5, 0, 0) FANOUT_363 (N3942, {N3942_0, N3942_1, N3942_2, N3942_3, N3942_4});
fanout_n #(7, 0, 0) FANOUT_364 (N3948, {N3948_0, N3948_1, N3948_2, N3948_3, N3948_4, N3948_5, N3948_6});
fanout_n #(5, 0, 0) FANOUT_365 (N3956, {N3956_0, N3956_1, N3956_2, N3956_3, N3956_4});
fanout_n #(5, 0, 0) FANOUT_366 (N3962, {N3962_0, N3962_1, N3962_2, N3962_3, N3962_4});
fanout_n #(6, 0, 0) FANOUT_367 (N3968, {N3968_0, N3968_1, N3968_2, N3968_3, N3968_4, N3968_5});
fanout_n #(2, 0, 0) FANOUT_368 (N3984, {N3984_0, N3984_1});
fanout_n #(2, 0, 0) FANOUT_369 (N4008, {N4008_0, N4008_1});
fanout_n #(2, 0, 0) FANOUT_370 (N4011, {N4011_0, N4011_1});
fanout_n #(2, 0, 0) FANOUT_371 (N4021, {N4021_0, N4021_1});
fanout_n #(2, 0, 0) FANOUT_372 (N4067, {N4067_0, N4067_1});
fanout_n #(3, 0, 0) FANOUT_373 (N4080, {N4080_0, N4080_1, N4080_2});
fanout_n #(2, 0, 0) FANOUT_374 (N4088, {N4088_0, N4088_1});
fanout_n #(2, 0, 0) FANOUT_375 (N4091, {N4091_0, N4091_1});
fanout_n #(2, 0, 0) FANOUT_376 (N4094, {N4094_0, N4094_1});
fanout_n #(2, 0, 0) FANOUT_377 (N4097, {N4097_0, N4097_1});
fanout_n #(2, 0, 0) FANOUT_378 (N4100, {N4100_0, N4100_1});
fanout_n #(2, 0, 0) FANOUT_379 (N4103, {N4103_0, N4103_1});
fanout_n #(2, 0, 0) FANOUT_380 (N4106, {N4106_0, N4106_1});
fanout_n #(2, 0, 0) FANOUT_381 (N4109, {N4109_0, N4109_1});
fanout_n #(2, 0, 0) FANOUT_382 (N4144, {N4144_0, N4144_1});
fanout_n #(2, 0, 0) FANOUT_383 (N4147, {N4147_0, N4147_1});
fanout_n #(2, 0, 0) FANOUT_384 (N4150, {N4150_0, N4150_1});
fanout_n #(2, 0, 0) FANOUT_385 (N4153, {N4153_0, N4153_1});
fanout_n #(2, 0, 0) FANOUT_386 (N4156, {N4156_0, N4156_1});
fanout_n #(2, 0, 0) FANOUT_387 (N4159, {N4159_0, N4159_1});
fanout_n #(2, 0, 0) FANOUT_388 (N4188, {N4188_0, N4188_1});
fanout_n #(2, 0, 0) FANOUT_389 (N4191, {N4191_0, N4191_1});
fanout_n #(2, 0, 0) FANOUT_390 (N4200, {N4200_0, N4200_1});
fanout_n #(2, 0, 0) FANOUT_391 (N4203, {N4203_0, N4203_1});
fanout_n #(2, 0, 0) FANOUT_392 (N4206, {N4206_0, N4206_1});
fanout_n #(2, 0, 0) FANOUT_393 (N4209, {N4209_0, N4209_1});
fanout_n #(2, 0, 0) FANOUT_394 (N4212, {N4212_0, N4212_1});
fanout_n #(2, 0, 0) FANOUT_395 (N4215, {N4215_0, N4215_1});
fanout_n #(2, 0, 0) FANOUT_396 (N4219, {N4219_0, N4219_1});
fanout_n #(2, 0, 0) FANOUT_397 (N4225, {N4225_0, N4225_1});
fanout_n #(2, 0, 0) FANOUT_398 (N4228, {N4228_0, N4228_1});
fanout_n #(2, 0, 0) FANOUT_399 (N4231, {N4231_0, N4231_1});
fanout_n #(2, 0, 0) FANOUT_400 (N4234, {N4234_0, N4234_1});
fanout_n #(2, 0, 0) FANOUT_401 (N4237, {N4237_0, N4237_1});
fanout_n #(2, 0, 0) FANOUT_402 (N4240, {N4240_0, N4240_1});
fanout_n #(2, 0, 0) FANOUT_403 (N4243, {N4243_0, N4243_1});
fanout_n #(2, 0, 0) FANOUT_404 (N4246, {N4246_0, N4246_1});
fanout_n #(2, 0, 0) FANOUT_405 (N4249, {N4249_0, N4249_1});
fanout_n #(2, 0, 0) FANOUT_406 (N4252, {N4252_0, N4252_1});
fanout_n #(2, 0, 0) FANOUT_407 (N4255, {N4255_0, N4255_1});
fanout_n #(2, 0, 0) FANOUT_408 (N4258, {N4258_0, N4258_1});
fanout_n #(2, 0, 0) FANOUT_409 (N4264, {N4264_0, N4264_1});
fanout_n #(3, 0, 0) FANOUT_410 (N4280, {N4280_0, N4280_1, N4280_2});
fanout_n #(5, 0, 0) FANOUT_411 (N4284, {N4284_0, N4284_1, N4284_2, N4284_3, N4284_4});
fanout_n #(6, 0, 0) FANOUT_412 (N4290, {N4290_0, N4290_1, N4290_2, N4290_3, N4290_4, N4290_5});
fanout_n #(2, 0, 0) FANOUT_413 (N4298, {N4298_0, N4298_1});
fanout_n #(3, 0, 0) FANOUT_414 (N4301, {N4301_0, N4301_1, N4301_2});
fanout_n #(4, 0, 0) FANOUT_415 (N4305, {N4305_0, N4305_1, N4305_2, N4305_3});
fanout_n #(5, 0, 0) FANOUT_416 (N4310, {N4310_0, N4310_1, N4310_2, N4310_3, N4310_4});
fanout_n #(3, 0, 0) FANOUT_417 (N4316, {N4316_0, N4316_1, N4316_2});
fanout_n #(4, 0, 0) FANOUT_418 (N4320, {N4320_0, N4320_1, N4320_2, N4320_3});
fanout_n #(5, 0, 0) FANOUT_419 (N4325, {N4325_0, N4325_1, N4325_2, N4325_3, N4325_4});
fanout_n #(3, 0, 0) FANOUT_420 (N4332, {N4332_0, N4332_1, N4332_2});
fanout_n #(5, 0, 0) FANOUT_421 (N4336, {N4336_0, N4336_1, N4336_2, N4336_3, N4336_4});
fanout_n #(6, 0, 0) FANOUT_422 (N4342, {N4342_0, N4342_1, N4342_2, N4342_3, N4342_4, N4342_5});
fanout_n #(7, 0, 0) FANOUT_423 (N4349, {N4349_0, N4349_1, N4349_2, N4349_3, N4349_4, N4349_5, N4349_6});
fanout_n #(6, 0, 0) FANOUT_424 (N4357, {N4357_0, N4357_1, N4357_2, N4357_3, N4357_4, N4357_5});
fanout_n #(10, 0, 0) FANOUT_425 (N4364, {N4364_0, N4364_1, N4364_2, N4364_3, N4364_4, N4364_5, N4364_6, N4364_7, N4364_8, N4364_9});
fanout_n #(3, 0, 0) FANOUT_426 (N4375, {N4375_0, N4375_1, N4375_2});
fanout_n #(5, 0, 0) FANOUT_427 (N4379, {N4379_0, N4379_1, N4379_2, N4379_3, N4379_4});
fanout_n #(6, 0, 0) FANOUT_428 (N4385, {N4385_0, N4385_1, N4385_2, N4385_3, N4385_4, N4385_5});
fanout_n #(3, 0, 0) FANOUT_429 (N4396, {N4396_0, N4396_1, N4396_2});
fanout_n #(4, 0, 0) FANOUT_430 (N4400, {N4400_0, N4400_1, N4400_2, N4400_3});
fanout_n #(6, 0, 0) FANOUT_431 (N4405, {N4405_0, N4405_1, N4405_2, N4405_3, N4405_4, N4405_5});
fanout_n #(5, 0, 0) FANOUT_432 (N4412, {N4412_0, N4412_1, N4412_2, N4412_3, N4412_4});
fanout_n #(6, 0, 0) FANOUT_433 (N4418, {N4418_0, N4418_1, N4418_2, N4418_3, N4418_4, N4418_5});
fanout_n #(10, 0, 0) FANOUT_434 (N4425, {N4425_0, N4425_1, N4425_2, N4425_3, N4425_4, N4425_5, N4425_6, N4425_7, N4425_8, N4425_9});
fanout_n #(3, 0, 0) FANOUT_435 (N4436, {N4436_0, N4436_1, N4436_2});
fanout_n #(4, 0, 0) FANOUT_436 (N4440, {N4440_0, N4440_1, N4440_2, N4440_3});
fanout_n #(5, 0, 0) FANOUT_437 (N4445, {N4445_0, N4445_1, N4445_2, N4445_3, N4445_4});
fanout_n #(5, 0, 0) FANOUT_438 (N4456, {N4456_0, N4456_1, N4456_2, N4456_3, N4456_4});
fanout_n #(6, 0, 0) FANOUT_439 (N4462, {N4462_0, N4462_1, N4462_2, N4462_3, N4462_4, N4462_5});
fanout_n #(7, 0, 0) FANOUT_440 (N4469, {N4469_0, N4469_1, N4469_2, N4469_3, N4469_4, N4469_5, N4469_6});
fanout_n #(6, 0, 0) FANOUT_441 (N4477, {N4477_0, N4477_1, N4477_2, N4477_3, N4477_4, N4477_5});
fanout_n #(2, 0, 0) FANOUT_442 (N4512, {N4512_0, N4512_1});
fanout_n #(3, 0, 0) FANOUT_443 (N4524, {N4524_0, N4524_1, N4524_2});
fanout_n #(3, 0, 0) FANOUT_444 (N4532, {N4532_0, N4532_1, N4532_2});
fanout_n #(2, 0, 0) FANOUT_445 (N4548, {N4548_0, N4548_1});
fanout_n #(2, 0, 0) FANOUT_446 (N4551, {N4551_0, N4551_1});
fanout_n #(2, 0, 0) FANOUT_447 (N4554, {N4554_0, N4554_1});
fanout_n #(2, 0, 0) FANOUT_448 (N4557, {N4557_0, N4557_1});
fanout_n #(2, 0, 0) FANOUT_449 (N4560, {N4560_0, N4560_1});
fanout_n #(2, 0, 0) FANOUT_450 (N4563, {N4563_0, N4563_1});
fanout_n #(2, 0, 0) FANOUT_451 (N4566, {N4566_0, N4566_1});
fanout_n #(2, 0, 0) FANOUT_452 (N4569, {N4569_0, N4569_1});
fanout_n #(2, 0, 0) FANOUT_453 (N4572, {N4572_0, N4572_1});
fanout_n #(2, 0, 0) FANOUT_454 (N4575, {N4575_0, N4575_1});
fanout_n #(2, 0, 0) FANOUT_455 (N4578, {N4578_0, N4578_1});
fanout_n #(2, 0, 0) FANOUT_456 (N4581, {N4581_0, N4581_1});
fanout_n #(2, 0, 0) FANOUT_457 (N4584, {N4584_0, N4584_1});
fanout_n #(2, 0, 0) FANOUT_458 (N4587, {N4587_0, N4587_1});
fanout_n #(2, 0, 0) FANOUT_459 (N4590, {N4590_0, N4590_1});
fanout_n #(2, 0, 0) FANOUT_460 (N4593, {N4593_0, N4593_1});
fanout_n #(2, 0, 0) FANOUT_461 (N4596, {N4596_0, N4596_1});
fanout_n #(2, 0, 0) FANOUT_462 (N4599, {N4599_0, N4599_1});
fanout_n #(2, 0, 0) FANOUT_463 (N4602, {N4602_0, N4602_1});
fanout_n #(2, 0, 0) FANOUT_464 (N4605, {N4605_0, N4605_1});
fanout_n #(2, 0, 0) FANOUT_465 (N4608, {N4608_0, N4608_1});
fanout_n #(2, 0, 0) FANOUT_466 (N4611, {N4611_0, N4611_1});
fanout_n #(2, 0, 0) FANOUT_467 (N4614, {N4614_0, N4614_1});
fanout_n #(2, 0, 0) FANOUT_468 (N4617, {N4617_0, N4617_1});
fanout_n #(2, 0, 0) FANOUT_469 (N4621, {N4621_0, N4621_1});
fanout_n #(2, 0, 0) FANOUT_470 (N4624, {N4624_0, N4624_1});
fanout_n #(2, 0, 0) FANOUT_471 (N4627, {N4627_0, N4627_1});
fanout_n #(2, 0, 0) FANOUT_472 (N4630, {N4630_0, N4630_1});
fanout_n #(2, 0, 0) FANOUT_473 (N4633, {N4633_0, N4633_1});
fanout_n #(2, 0, 0) FANOUT_474 (N4637, {N4637_0, N4637_1});
fanout_n #(2, 0, 0) FANOUT_475 (N4640, {N4640_0, N4640_1});
fanout_n #(2, 0, 0) FANOUT_476 (N4643, {N4643_0, N4643_1});
fanout_n #(2, 0, 0) FANOUT_477 (N4646, {N4646_0, N4646_1});
fanout_n #(2, 0, 0) FANOUT_478 (N4649, {N4649_0, N4649_1});
fanout_n #(2, 0, 0) FANOUT_479 (N4652, {N4652_0, N4652_1});
fanout_n #(2, 0, 0) FANOUT_480 (N4655, {N4655_0, N4655_1});
fanout_n #(2, 0, 0) FANOUT_481 (N4658, {N4658_0, N4658_1});
fanout_n #(2, 0, 0) FANOUT_482 (N4662, {N4662_0, N4662_1});
fanout_n #(2, 0, 0) FANOUT_483 (N4665, {N4665_0, N4665_1});
fanout_n #(2, 0, 0) FANOUT_484 (N4668, {N4668_0, N4668_1});
fanout_n #(2, 0, 0) FANOUT_485 (N4671, {N4671_0, N4671_1});
fanout_n #(2, 0, 0) FANOUT_486 (N4674, {N4674_0, N4674_1});
fanout_n #(2, 0, 0) FANOUT_487 (N4677, {N4677_0, N4677_1});
fanout_n #(2, 0, 0) FANOUT_488 (N4680, {N4680_0, N4680_1});
fanout_n #(2, 0, 0) FANOUT_489 (N4683, {N4683_0, N4683_1});
fanout_n #(2, 0, 0) FANOUT_490 (N4686, {N4686_0, N4686_1});
fanout_n #(2, 0, 0) FANOUT_491 (N4689, {N4689_0, N4689_1});
fanout_n #(2, 0, 0) FANOUT_492 (N4692, {N4692_0, N4692_1});
fanout_n #(2, 0, 0) FANOUT_493 (N4695, {N4695_0, N4695_1});
fanout_n #(2, 0, 0) FANOUT_494 (N4698, {N4698_0, N4698_1});
fanout_n #(2, 0, 0) FANOUT_495 (N4939, {N4939_0, N4939_1});
fanout_n #(2, 0, 0) FANOUT_496 (N5049, {N5049_0, N5049_1});
fanout_n #(2, 0, 0) FANOUT_497 (N5150, {N5150_0, N5150_1});
fanout_n #(2, 0, 0) FANOUT_498 (N5157, {N5157_0, N5157_1});
fanout_n #(2, 0, 0) FANOUT_499 (N5166, {N5166_0, N5166_1});
fanout_n #(2, 0, 0) FANOUT_500 (N5169, {N5169_0, N5169_1});
fanout_n #(2, 0, 0) FANOUT_501 (N5173, {N5173_0, N5173_1});
fanout_n #(2, 0, 0) FANOUT_502 (N5177, {N5177_0, N5177_1});
fanout_n #(2, 0, 0) FANOUT_503 (N5180, {N5180_0, N5180_1});
fanout_n #(2, 0, 0) FANOUT_504 (N5183, {N5183_0, N5183_1});
fanout_n #(2, 0, 0) FANOUT_505 (N5186, {N5186_0, N5186_1});
fanout_n #(2, 0, 0) FANOUT_506 (N5189, {N5189_0, N5189_1});
fanout_n #(2, 0, 0) FANOUT_507 (N5192, {N5192_0, N5192_1});
fanout_n #(2, 0, 0) FANOUT_508 (N5195, {N5195_0, N5195_1});
fanout_n #(2, 0, 0) FANOUT_509 (N5199, {N5199_0, N5199_1});
fanout_n #(2, 0, 0) FANOUT_510 (N5202, {N5202_0, N5202_1});
fanout_n #(2, 0, 0) FANOUT_511 (N5205, {N5205_0, N5205_1});
fanout_n #(2, 0, 0) FANOUT_512 (N5208, {N5208_0, N5208_1});
fanout_n #(2, 0, 0) FANOUT_513 (N5211, {N5211_0, N5211_1});
fanout_n #(2, 0, 0) FANOUT_514 (N5214, {N5214_0, N5214_1});
fanout_n #(2, 0, 0) FANOUT_515 (N5217, {N5217_0, N5217_1});
fanout_n #(2, 0, 0) FANOUT_516 (N5220, {N5220_0, N5220_1});
fanout_n #(2, 0, 0) FANOUT_517 (N5236, {N5236_0, N5236_1});
fanout_n #(9, 0, 0) FANOUT_518 (N5264, {N5264_0, N5264_1, N5264_2, N5264_3, N5264_4, N5264_5, N5264_6, N5264_7, N5264_8});
fanout_n #(13, 0, 0) FANOUT_519 (N5284, {N5284_0, N5284_1, N5284_2, N5284_3, N5284_4, N5284_5, N5284_6, N5284_7, N5284_8, N5284_9, N5284_10, N5284_11, N5284_12});
fanout_n #(3, 0, 0) FANOUT_520 (N5315, {N5315_0, N5315_1, N5315_2});
fanout_n #(2, 0, 0) FANOUT_521 (N5319, {N5319_0, N5319_1});
fanout_n #(3, 0, 0) FANOUT_522 (N5324, {N5324_0, N5324_1, N5324_2});
fanout_n #(2, 0, 0) FANOUT_523 (N5328, {N5328_0, N5328_1});
fanout_n #(2, 0, 0) FANOUT_524 (N5346, {N5346_0, N5346_1});
fanout_n #(2, 0, 0) FANOUT_525 (N5371, {N5371_0, N5371_1});
fanout_n #(2, 0, 0) FANOUT_526 (N5374, {N5374_0, N5374_1});
fanout_n #(2, 0, 0) FANOUT_527 (N5377, {N5377_0, N5377_1});
fanout_n #(2, 0, 0) FANOUT_528 (N5382, {N5382_0, N5382_1});
fanout_n #(2, 0, 0) FANOUT_529 (N5385, {N5385_0, N5385_1});
fanout_n #(6, 0, 0) FANOUT_530 (N5389, {N5389_0, N5389_1, N5389_2, N5389_3, N5389_4, N5389_5});
fanout_n #(10, 0, 0) FANOUT_531 (N5396, {N5396_0, N5396_1, N5396_2, N5396_3, N5396_4, N5396_5, N5396_6, N5396_7, N5396_8, N5396_9});
fanout_n #(10, 0, 0) FANOUT_532 (N5407, {N5407_0, N5407_1, N5407_2, N5407_3, N5407_4, N5407_5, N5407_6, N5407_7, N5407_8, N5407_9});
fanout_n #(5, 0, 0) FANOUT_533 (N5418, {N5418_0, N5418_1, N5418_2, N5418_3, N5418_4});
fanout_n #(6, 0, 0) FANOUT_534 (N5424, {N5424_0, N5424_1, N5424_2, N5424_3, N5424_4, N5424_5});
fanout_n #(9, 0, 0) FANOUT_535 (N5431, {N5431_0, N5431_1, N5431_2, N5431_3, N5431_4, N5431_5, N5431_6, N5431_7, N5431_8});
fanout_n #(10, 0, 0) FANOUT_536 (N5441, {N5441_0, N5441_1, N5441_2, N5441_3, N5441_4, N5441_5, N5441_6, N5441_7, N5441_8, N5441_9});
fanout_n #(9, 0, 0) FANOUT_537 (N5452, {N5452_0, N5452_1, N5452_2, N5452_3, N5452_4, N5452_5, N5452_6, N5452_7, N5452_8});
fanout_n #(6, 0, 0) FANOUT_538 (N5462, {N5462_0, N5462_1, N5462_2, N5462_3, N5462_4, N5462_5});
fanout_n #(6, 0, 0) FANOUT_539 (N5470, {N5470_0, N5470_1, N5470_2, N5470_3, N5470_4, N5470_5});
fanout_n #(10, 0, 0) FANOUT_540 (N5477, {N5477_0, N5477_1, N5477_2, N5477_3, N5477_4, N5477_5, N5477_6, N5477_7, N5477_8, N5477_9});
fanout_n #(9, 0, 0) FANOUT_541 (N5488, {N5488_0, N5488_1, N5488_2, N5488_3, N5488_4, N5488_5, N5488_6, N5488_7, N5488_8});
fanout_n #(7, 0, 0) FANOUT_542 (N5498, {N5498_0, N5498_1, N5498_2, N5498_3, N5498_4, N5498_5, N5498_6});
fanout_n #(13, 0, 0) FANOUT_543 (N5506, {N5506_0, N5506_1, N5506_2, N5506_3, N5506_4, N5506_5, N5506_6, N5506_7, N5506_8, N5506_9, N5506_10, N5506_11, N5506_12});
fanout_n #(15, 0, 0) FANOUT_544 (N5520, {N5520_0, N5520_1, N5520_2, N5520_3, N5520_4, N5520_5, N5520_6, N5520_7, N5520_8, N5520_9, N5520_10, N5520_11, N5520_12, N5520_13, N5520_14});
fanout_n #(12, 0, 0) FANOUT_545 (N5536, {N5536_0, N5536_1, N5536_2, N5536_3, N5536_4, N5536_5, N5536_6, N5536_7, N5536_8, N5536_9, N5536_10, N5536_11});
fanout_n #(5, 0, 0) FANOUT_546 (N5549, {N5549_0, N5549_1, N5549_2, N5549_3, N5549_4});
fanout_n #(6, 0, 0) FANOUT_547 (N5555, {N5555_0, N5555_1, N5555_2, N5555_3, N5555_4, N5555_5});
fanout_n #(10, 0, 0) FANOUT_548 (N5562, {N5562_0, N5562_1, N5562_2, N5562_3, N5562_4, N5562_5, N5562_6, N5562_7, N5562_8, N5562_9});
fanout_n #(5, 0, 0) FANOUT_549 (N5573, {N5573_0, N5573_1, N5573_2, N5573_3, N5573_4});
fanout_n #(6, 0, 0) FANOUT_550 (N5579, {N5579_0, N5579_1, N5579_2, N5579_3, N5579_4, N5579_5});
fanout_n #(10, 0, 0) FANOUT_551 (N5595, {N5595_0, N5595_1, N5595_2, N5595_3, N5595_4, N5595_5, N5595_6, N5595_7, N5595_8, N5595_9});
fanout_n #(9, 0, 0) FANOUT_552 (N5606, {N5606_0, N5606_1, N5606_2, N5606_3, N5606_4, N5606_5, N5606_6, N5606_7, N5606_8});
fanout_n #(9, 0, 0) FANOUT_553 (N5624, {N5624_0, N5624_1, N5624_2, N5624_3, N5624_4, N5624_5, N5624_6, N5624_7, N5624_8});
fanout_n #(7, 0, 0) FANOUT_554 (N5634, {N5634_0, N5634_1, N5634_2, N5634_3, N5634_4, N5634_5, N5634_6});
fanout_n #(15, 0, 0) FANOUT_555 (N5655, {N5655_0, N5655_1, N5655_2, N5655_3, N5655_4, N5655_5, N5655_6, N5655_7, N5655_8, N5655_9, N5655_10, N5655_11, N5655_12, N5655_13, N5655_14});
fanout_n #(12, 0, 0) FANOUT_556 (N5671, {N5671_0, N5671_1, N5671_2, N5671_3, N5671_4, N5671_5, N5671_6, N5671_7, N5671_8, N5671_9, N5671_10, N5671_11});
fanout_n #(5, 0, 0) FANOUT_557 (N5684, {N5684_0, N5684_1, N5684_2, N5684_3, N5684_4});
fanout_n #(3, 0, 0) FANOUT_558 (N5692, {N5692_0, N5692_1, N5692_2});
fanout_n #(3, 0, 0) FANOUT_559 (N5696, {N5696_0, N5696_1, N5696_2});
fanout_n #(2, 0, 0) FANOUT_560 (N5700, {N5700_0, N5700_1});
fanout_n #(3, 0, 0) FANOUT_561 (N5703, {N5703_0, N5703_1, N5703_2});
fanout_n #(3, 0, 0) FANOUT_562 (N5707, {N5707_0, N5707_1, N5707_2});
fanout_n #(2, 0, 0) FANOUT_563 (N5711, {N5711_0, N5711_1});
fanout_n #(2, 0, 0) FANOUT_564 (N5736, {N5736_0, N5736_1});
fanout_n #(2, 0, 0) FANOUT_565 (N5739, {N5739_0, N5739_1});
fanout_n #(2, 0, 0) FANOUT_566 (N5742, {N5742_0, N5742_1});
fanout_n #(2, 0, 0) FANOUT_567 (N5745, {N5745_0, N5745_1});
fanout_n #(2, 0, 0) FANOUT_568 (N5756, {N5756_0, N5756_1});
fanout_n #(2, 0, 0) FANOUT_569 (N6025, {N6025_0, N6025_1});
fanout_n #(2, 0, 0) FANOUT_570 (N6028, {N6028_0, N6028_1});
fanout_n #(2, 0, 0) FANOUT_571 (N6031, {N6031_0, N6031_1});
fanout_n #(2, 0, 0) FANOUT_572 (N6034, {N6034_0, N6034_1});
fanout_n #(2, 0, 0) FANOUT_573 (N6037, {N6037_0, N6037_1});
fanout_n #(2, 0, 0) FANOUT_574 (N6040, {N6040_0, N6040_1});
fanout_n #(2, 0, 0) FANOUT_575 (N6045, {N6045_0, N6045_1});
fanout_n #(2, 0, 0) FANOUT_576 (N6048, {N6048_0, N6048_1});
fanout_n #(2, 0, 0) FANOUT_577 (N6051, {N6051_0, N6051_1});
fanout_n #(2, 0, 0) FANOUT_578 (N6054, {N6054_0, N6054_1});
fanout_n #(2, 0, 0) FANOUT_579 (N6080, {N6080_0, N6080_1});
fanout_n #(2, 0, 0) FANOUT_580 (N6091, {N6091_0, N6091_1});
fanout_n #(2, 0, 0) FANOUT_581 (N6108, {N6108_0, N6108_1});
fanout_n #(2, 0, 0) FANOUT_582 (N6117, {N6117_0, N6117_1});
fanout_n #(2, 0, 0) FANOUT_583 (N6140, {N6140_0, N6140_1});
fanout_n #(2, 0, 0) FANOUT_584 (N6149, {N6149_0, N6149_1});
fanout_n #(2, 0, 0) FANOUT_585 (N6164, {N6164_0, N6164_1});
fanout_n #(2, 0, 0) FANOUT_586 (N6168, {N6168_0, N6168_1});
fanout_n #(2, 0, 0) FANOUT_587 (N6175, {N6175_0, N6175_1});
fanout_n #(2, 0, 0) FANOUT_588 (N6197, {N6197_0, N6197_1});
fanout_n #(2, 0, 0) FANOUT_589 (N6200, {N6200_0, N6200_1});
fanout_n #(2, 0, 0) FANOUT_590 (N6203, {N6203_0, N6203_1});
fanout_n #(2, 0, 0) FANOUT_591 (N6206, {N6206_0, N6206_1});
fanout_n #(2, 0, 0) FANOUT_592 (N6209, {N6209_0, N6209_1});
fanout_n #(2, 0, 0) FANOUT_593 (N6212, {N6212_0, N6212_1});
fanout_n #(2, 0, 0) FANOUT_594 (N6215, {N6215_0, N6215_1});
fanout_n #(2, 0, 0) FANOUT_595 (N6218, {N6218_0, N6218_1});
fanout_n #(2, 0, 0) FANOUT_596 (N6238, {N6238_0, N6238_1});
fanout_n #(2, 0, 0) FANOUT_597 (N6241, {N6241_0, N6241_1});
fanout_n #(2, 0, 0) FANOUT_598 (N6244, {N6244_0, N6244_1});
fanout_n #(2, 0, 0) FANOUT_599 (N6247, {N6247_0, N6247_1});
fanout_n #(2, 0, 0) FANOUT_600 (N6250, {N6250_0, N6250_1});
fanout_n #(2, 0, 0) FANOUT_601 (N6253, {N6253_0, N6253_1});
fanout_n #(2, 0, 0) FANOUT_602 (N6256, {N6256_0, N6256_1});
fanout_n #(2, 0, 0) FANOUT_603 (N6259, {N6259_0, N6259_1});
fanout_n #(2, 0, 0) FANOUT_604 (N6262, {N6262_0, N6262_1});
fanout_n #(2, 0, 0) FANOUT_605 (N6265, {N6265_0, N6265_1});
fanout_n #(2, 0, 0) FANOUT_606 (N6268, {N6268_0, N6268_1});
fanout_n #(2, 0, 0) FANOUT_607 (N6271, {N6271_0, N6271_1});
fanout_n #(2, 0, 0) FANOUT_608 (N6274, {N6274_0, N6274_1});
fanout_n #(2, 0, 0) FANOUT_609 (N6277, {N6277_0, N6277_1});
fanout_n #(2, 0, 0) FANOUT_610 (N6280, {N6280_0, N6280_1});
fanout_n #(2, 0, 0) FANOUT_611 (N6283, {N6283_0, N6283_1});
fanout_n #(2, 0, 0) FANOUT_612 (N6286, {N6286_0, N6286_1});
fanout_n #(2, 0, 0) FANOUT_613 (N6289, {N6289_0, N6289_1});
fanout_n #(2, 0, 0) FANOUT_614 (N6292, {N6292_0, N6292_1});
fanout_n #(2, 0, 0) FANOUT_615 (N6295, {N6295_0, N6295_1});
fanout_n #(2, 0, 0) FANOUT_616 (N6298, {N6298_0, N6298_1});
fanout_n #(2, 0, 0) FANOUT_617 (N6301, {N6301_0, N6301_1});
fanout_n #(2, 0, 0) FANOUT_618 (N6304, {N6304_0, N6304_1});
fanout_n #(2, 0, 0) FANOUT_619 (N6307, {N6307_0, N6307_1});
fanout_n #(2, 0, 0) FANOUT_620 (N6310, {N6310_0, N6310_1});
fanout_n #(2, 0, 0) FANOUT_621 (N6313, {N6313_0, N6313_1});
fanout_n #(2, 0, 0) FANOUT_622 (N6316, {N6316_0, N6316_1});
fanout_n #(2, 0, 0) FANOUT_623 (N6319, {N6319_0, N6319_1});
fanout_n #(2, 0, 0) FANOUT_624 (N6322, {N6322_0, N6322_1});
fanout_n #(2, 0, 0) FANOUT_625 (N6325, {N6325_0, N6325_1});
fanout_n #(2, 0, 0) FANOUT_626 (N6328, {N6328_0, N6328_1});
fanout_n #(2, 0, 0) FANOUT_627 (N6331, {N6331_0, N6331_1});
fanout_n #(2, 0, 0) FANOUT_628 (N6335, {N6335_0, N6335_1});
fanout_n #(2, 0, 0) FANOUT_629 (N6338, {N6338_0, N6338_1});
fanout_n #(2, 0, 0) FANOUT_630 (N6341, {N6341_0, N6341_1});
fanout_n #(2, 0, 0) FANOUT_631 (N6344, {N6344_0, N6344_1});
fanout_n #(2, 0, 0) FANOUT_632 (N6347, {N6347_0, N6347_1});
fanout_n #(2, 0, 0) FANOUT_633 (N6350, {N6350_0, N6350_1});
fanout_n #(2, 0, 0) FANOUT_634 (N6353, {N6353_0, N6353_1});
fanout_n #(2, 0, 0) FANOUT_635 (N6356, {N6356_0, N6356_1});
fanout_n #(2, 0, 0) FANOUT_636 (N6359, {N6359_0, N6359_1});
fanout_n #(2, 0, 0) FANOUT_637 (N6364, {N6364_0, N6364_1});
fanout_n #(2, 0, 0) FANOUT_638 (N6367, {N6367_0, N6367_1});
fanout_n #(2, 0, 0) FANOUT_639 (N6370, {N6370_0, N6370_1});
fanout_n #(2, 0, 0) FANOUT_640 (N6397, {N6397_0, N6397_1});
fanout_n #(2, 0, 0) FANOUT_641 (N6411, {N6411_0, N6411_1});
fanout_n #(3, 0, 0) FANOUT_642 (N6415, {N6415_0, N6415_1, N6415_2});
fanout_n #(2, 0, 0) FANOUT_643 (N6419, {N6419_0, N6419_1});
fanout_n #(2, 0, 0) FANOUT_644 (N6427, {N6427_0, N6427_1});
fanout_n #(2, 0, 0) FANOUT_645 (N6437, {N6437_0, N6437_1});
fanout_n #(3, 0, 0) FANOUT_646 (N6441, {N6441_0, N6441_1, N6441_2});
fanout_n #(2, 0, 0) FANOUT_647 (N6445, {N6445_0, N6445_1});
fanout_n #(2, 0, 0) FANOUT_648 (N6466, {N6466_0, N6466_1});
fanout_n #(2, 0, 0) FANOUT_649 (N6478, {N6478_0, N6478_1});
fanout_n #(2, 0, 0) FANOUT_650 (N6482, {N6482_0, N6482_1});
fanout_n #(2, 0, 0) FANOUT_651 (N6486, {N6486_0, N6486_1});
fanout_n #(2, 0, 0) FANOUT_652 (N6490, {N6490_0, N6490_1});
fanout_n #(2, 0, 0) FANOUT_653 (N6494, {N6494_0, N6494_1});
fanout_n #(2, 0, 0) FANOUT_654 (N6500, {N6500_0, N6500_1});
fanout_n #(2, 0, 0) FANOUT_655 (N6504, {N6504_0, N6504_1});
fanout_n #(2, 0, 0) FANOUT_656 (N6508, {N6508_0, N6508_1});
fanout_n #(2, 0, 0) FANOUT_657 (N6512, {N6512_0, N6512_1});
fanout_n #(2, 0, 0) FANOUT_658 (N6516, {N6516_0, N6516_1});
fanout_n #(2, 0, 0) FANOUT_659 (N6526, {N6526_0, N6526_1});
fanout_n #(2, 0, 0) FANOUT_660 (N6536, {N6536_0, N6536_1});
fanout_n #(2, 0, 0) FANOUT_661 (N6539, {N6539_0, N6539_1});
fanout_n #(2, 0, 0) FANOUT_662 (N6553, {N6553_0, N6553_1});
fanout_n #(2, 0, 0) FANOUT_663 (N6556, {N6556_0, N6556_1});
fanout_n #(2, 0, 0) FANOUT_664 (N6566, {N6566_0, N6566_1});
fanout_n #(2, 0, 0) FANOUT_665 (N6569, {N6569_0, N6569_1});
fanout_n #(2, 0, 0) FANOUT_666 (N6572, {N6572_0, N6572_1});
fanout_n #(2, 0, 0) FANOUT_667 (N6575, {N6575_0, N6575_1});
fanout_n #(2, 0, 0) FANOUT_668 (N6580, {N6580_0, N6580_1});
fanout_n #(2, 0, 0) FANOUT_669 (N6584, {N6584_0, N6584_1});
fanout_n #(2, 0, 0) FANOUT_670 (N6587, {N6587_0, N6587_1});
fanout_n #(2, 0, 0) FANOUT_671 (N6592, {N6592_0, N6592_1});
fanout_n #(2, 0, 0) FANOUT_672 (N6599, {N6599_0, N6599_1});
fanout_n #(2, 0, 0) FANOUT_673 (N6606, {N6606_0, N6606_1});
fanout_n #(2, 0, 0) FANOUT_674 (N6609, {N6609_0, N6609_1});
fanout_n #(2, 0, 0) FANOUT_675 (N6619, {N6619_0, N6619_1});
fanout_n #(2, 0, 0) FANOUT_676 (N6622, {N6622_0, N6622_1});
fanout_n #(2, 0, 0) FANOUT_677 (N6634, {N6634_0, N6634_1});
fanout_n #(2, 0, 0) FANOUT_678 (N6637, {N6637_0, N6637_1});
fanout_n #(2, 0, 0) FANOUT_679 (N6724, {N6724_0, N6724_1});
fanout_n #(2, 0, 0) FANOUT_680 (N6792, {N6792_0, N6792_1});
fanout_n #(2, 0, 0) FANOUT_681 (N6795, {N6795_0, N6795_1});
fanout_n #(5, 0, 0) FANOUT_682 (N6817, {N6817_0, N6817_1, N6817_2, N6817_3, N6817_4});
fanout_n #(2, 0, 0) FANOUT_683 (N6831, {N6831_0, N6831_1});
fanout_n #(5, 0, 0) FANOUT_684 (N6844, {N6844_0, N6844_1, N6844_2, N6844_3, N6844_4});
fanout_n #(2, 0, 0) FANOUT_685 (N6857, {N6857_0, N6857_1});
fanout_n #(5, 0, 0) FANOUT_686 (N6866, {N6866_0, N6866_1, N6866_2, N6866_3, N6866_4});
fanout_n #(2, 0, 0) FANOUT_687 (N6881, {N6881_0, N6881_1});
fanout_n #(2, 0, 0) FANOUT_688 (N6885, {N6885_0, N6885_1});
fanout_n #(2, 0, 0) FANOUT_689 (N6891, {N6891_0, N6891_1});
fanout_n #(2, 0, 0) FANOUT_690 (N6897, {N6897_0, N6897_1});
fanout_n #(2, 0, 0) FANOUT_691 (N6901, {N6901_0, N6901_1});
fanout_n #(2, 0, 0) FANOUT_692 (N6905, {N6905_0, N6905_1});
fanout_n #(2, 0, 0) FANOUT_693 (N6909, {N6909_0, N6909_1});
fanout_n #(2, 0, 0) FANOUT_694 (N6916, {N6916_0, N6916_1});
fanout_n #(2, 0, 0) FANOUT_695 (N6932, {N6932_0, N6932_1});
fanout_n #(2, 0, 0) FANOUT_696 (N6967, {N6967_0, N6967_1});
fanout_n #(3, 0, 0) FANOUT_697 (N6979, {N6979_0, N6979_1, N6979_2});
fanout_n #(2, 0, 0) FANOUT_698 (N7003, {N7003_0, N7003_1});
fanout_n #(2, 0, 0) FANOUT_699 (N7006, {N7006_0, N7006_1});
fanout_n #(4, 0, 0) FANOUT_700 (N7023, {N7023_0, N7023_1, N7023_2, N7023_3});
fanout_n #(2, 0, 0) FANOUT_701 (N7028, {N7028_0, N7028_1});
fanout_n #(2, 0, 0) FANOUT_702 (N7031, {N7031_0, N7031_1});
fanout_n #(2, 0, 0) FANOUT_703 (N7034, {N7034_0, N7034_1});
fanout_n #(2, 0, 0) FANOUT_704 (N7037, {N7037_0, N7037_1});
fanout_n #(2, 0, 0) FANOUT_705 (N7041, {N7041_0, N7041_1});
fanout_n #(4, 0, 0) FANOUT_706 (N7049, {N7049_0, N7049_1, N7049_2, N7049_3});
fanout_n #(2, 0, 0) FANOUT_707 (N7054, {N7054_0, N7054_1});
fanout_n #(2, 0, 0) FANOUT_708 (N7057, {N7057_0, N7057_1});
fanout_n #(2, 0, 0) FANOUT_709 (N7060, {N7060_0, N7060_1});
fanout_n #(2, 0, 0) FANOUT_710 (N7065, {N7065_0, N7065_1});
fanout_n #(2, 0, 0) FANOUT_711 (N7076, {N7076_0, N7076_1});
fanout_n #(2, 0, 0) FANOUT_712 (N7080, {N7080_0, N7080_1});
fanout_n #(2, 0, 0) FANOUT_713 (N7090, {N7090_0, N7090_1});
fanout_n #(2, 0, 0) FANOUT_714 (N7094, {N7094_0, N7094_1});
fanout_n #(2, 0, 0) FANOUT_715 (N7097, {N7097_0, N7097_1});
fanout_n #(2, 0, 0) FANOUT_716 (N7101, {N7101_0, N7101_1});
fanout_n #(5, 0, 0) FANOUT_717 (N7190, {N7190_0, N7190_1, N7190_2, N7190_3, N7190_4});
fanout_n #(5, 0, 0) FANOUT_718 (N7198, {N7198_0, N7198_1, N7198_2, N7198_3, N7198_4});
fanout_n #(2, 0, 0) FANOUT_719 (N7209, {N7209_0, N7209_1});
fanout_n #(2, 0, 0) FANOUT_720 (N7212, {N7212_0, N7212_1});
fanout_n #(2, 0, 0) FANOUT_721 (N7219, {N7219_0, N7219_1});
fanout_n #(2, 0, 0) FANOUT_722 (N7222, {N7222_0, N7222_1});
fanout_n #(2, 0, 0) FANOUT_723 (N7225, {N7225_0, N7225_1});
fanout_n #(2, 0, 0) FANOUT_724 (N7236, {N7236_0, N7236_1});
fanout_n #(2, 0, 0) FANOUT_725 (N7239, {N7239_0, N7239_1});
fanout_n #(2, 0, 0) FANOUT_726 (N7242, {N7242_0, N7242_1});
fanout_n #(2, 0, 0) FANOUT_727 (N7245, {N7245_0, N7245_1});
fanout_n #(6, 0, 0) FANOUT_728 (N7250, {N7250_0, N7250_1, N7250_2, N7250_3, N7250_4, N7250_5});
fanout_n #(2, 0, 0) FANOUT_729 (N7257, {N7257_0, N7257_1});
fanout_n #(2, 0, 0) FANOUT_730 (N7260, {N7260_0, N7260_1});
fanout_n #(2, 0, 0) FANOUT_731 (N7263, {N7263_0, N7263_1});
fanout_n #(5, 0, 0) FANOUT_732 (N7270, {N7270_0, N7270_1, N7270_2, N7270_3, N7270_4});
fanout_n #(5, 0, 0) FANOUT_733 (N7276, {N7276_0, N7276_1, N7276_2, N7276_3, N7276_4});
fanout_n #(5, 0, 0) FANOUT_734 (N7282, {N7282_0, N7282_1, N7282_2, N7282_3, N7282_4});
fanout_n #(5, 0, 0) FANOUT_735 (N7288, {N7288_0, N7288_1, N7288_2, N7288_3, N7288_4});
fanout_n #(5, 0, 0) FANOUT_736 (N7294, {N7294_0, N7294_1, N7294_2, N7294_3, N7294_4});
fanout_n #(2, 0, 0) FANOUT_737 (N7301, {N7301_0, N7301_1});
fanout_n #(5, 0, 0) FANOUT_738 (N7304, {N7304_0, N7304_1, N7304_2, N7304_3, N7304_4});
fanout_n #(5, 0, 0) FANOUT_739 (N7310, {N7310_0, N7310_1, N7310_2, N7310_3, N7310_4});
fanout_n #(2, 0, 0) FANOUT_740 (N7394, {N7394_0, N7394_1});
fanout_n #(2, 0, 0) FANOUT_741 (N7397, {N7397_0, N7397_1});
fanout_n #(2, 0, 0) FANOUT_742 (N7402, {N7402_0, N7402_1});
fanout_n #(2, 0, 0) FANOUT_743 (N7409, {N7409_0, N7409_1});
fanout_n #(2, 0, 0) FANOUT_744 (N7412, {N7412_0, N7412_1});
fanout_n #(2, 0, 0) FANOUT_745 (N7421, {N7421_0, N7421_1});
fanout_n #(2, 0, 0) FANOUT_746 (N7489, {N7489_0, N7489_1});
fanout_n #(5, 0, 0) FANOUT_747 (N7531, {N7531_0, N7531_1, N7531_2, N7531_3, N7531_4});
fanout_n #(5, 0, 0) FANOUT_748 (N7537, {N7537_0, N7537_1, N7537_2, N7537_3, N7537_4});
fanout_n #(5, 0, 0) FANOUT_749 (N7543, {N7543_0, N7543_1, N7543_2, N7543_3, N7543_4});
fanout_n #(5, 0, 0) FANOUT_750 (N7549, {N7549_0, N7549_1, N7549_2, N7549_3, N7549_4});
fanout_n #(5, 0, 0) FANOUT_751 (N7555, {N7555_0, N7555_1, N7555_2, N7555_3, N7555_4});
fanout_n #(5, 0, 0) FANOUT_752 (N7561, {N7561_0, N7561_1, N7561_2, N7561_3, N7561_4});
fanout_n #(5, 0, 0) FANOUT_753 (N7567, {N7567_0, N7567_1, N7567_2, N7567_3, N7567_4});
fanout_n #(5, 0, 0) FANOUT_754 (N7573, {N7573_0, N7573_1, N7573_2, N7573_3, N7573_4});
fanout_n #(2, 0, 0) FANOUT_755 (N7579, {N7579_0, N7579_1});
fanout_n #(2, 0, 0) FANOUT_756 (N7582, {N7582_0, N7582_1});
fanout_n #(2, 0, 0) FANOUT_757 (N7589, {N7589_0, N7589_1});
fanout_n #(2, 0, 0) FANOUT_758 (N7592, {N7592_0, N7592_1});
fanout_n #(2, 0, 0) FANOUT_759 (N7595, {N7595_0, N7595_1});
fanout_n #(2, 0, 0) FANOUT_760 (N7712, {N7712_0, N7712_1});
fanout_n #(2, 0, 0) FANOUT_761 (N7715, {N7715_0, N7715_1});
fanout_n #(2, 0, 0) FANOUT_762 (N7724, {N7724_0, N7724_1});
fanout_n #(2, 0, 0) FANOUT_763 (N7762, {N7762_0, N7762_1});
fanout_n #(2, 0, 0) FANOUT_764 (N7765, {N7765_0, N7765_1});
fanout_n #(2, 0, 0) FANOUT_765 (N7772, {N7772_0, N7772_1});
fanout_n #(2, 0, 0) FANOUT_766 (N7775, {N7775_0, N7775_1});
fanout_n #(2, 0, 0) FANOUT_767 (N7778, {N7778_0, N7778_1});
fanout_n #(2, 0, 0) FANOUT_768 (N7800, {N7800_0, N7800_1});
fanout_n #(2, 0, 0) FANOUT_769 (N7803, {N7803_0, N7803_1});
fanout_n #(2, 0, 0) FANOUT_770 (N7812, {N7812_0, N7812_1});
fanout_n #(2, 0, 0) FANOUT_771 (N7826, {N7826_0, N7826_1});
fanout_n #(2, 0, 0) FANOUT_772 (N7829, {N7829_0, N7829_1});
fanout_n #(2, 0, 0) FANOUT_773 (N7836, {N7836_0, N7836_1});
fanout_n #(2, 0, 0) FANOUT_774 (N7839, {N7839_0, N7839_1});
fanout_n #(2, 0, 0) FANOUT_775 (N7842, {N7842_0, N7842_1});
fanout_n #(2, 0, 0) FANOUT_776 (N7864, {N7864_0, N7864_1});
fanout_n #(2, 0, 0) FANOUT_777 (N7867, {N7867_0, N7867_1});
fanout_n #(2, 0, 0) FANOUT_778 (N7876, {N7876_0, N7876_1});
fanout_n #(2, 0, 0) FANOUT_779 (N7890, {N7890_0, N7890_1});
fanout_n #(2, 0, 0) FANOUT_780 (N7893, {N7893_0, N7893_1});
fanout_n #(2, 0, 0) FANOUT_781 (N7900, {N7900_0, N7900_1});
fanout_n #(2, 0, 0) FANOUT_782 (N7903, {N7903_0, N7903_1});
fanout_n #(2, 0, 0) FANOUT_783 (N7906, {N7906_0, N7906_1});
fanout_n #(2, 0, 0) FANOUT_784 (N7932, {N7932_0, N7932_1});
fanout_n #(2, 0, 0) FANOUT_785 (N7935, {N7935_0, N7935_1});
fanout_n #(2, 0, 0) FANOUT_786 (N7940, {N7940_0, N7940_1});
fanout_n #(2, 0, 0) FANOUT_787 (N7954, {N7954_0, N7954_1});
fanout_n #(2, 0, 0) FANOUT_788 (N7957, {N7957_0, N7957_1});
fanout_n #(2, 0, 0) FANOUT_789 (N7960, {N7960_0, N7960_1});
fanout_n #(2, 0, 0) FANOUT_790 (N7963, {N7963_0, N7963_1});
fanout_n #(2, 0, 0) FANOUT_791 (N7970, {N7970_0, N7970_1});
fanout_n #(2, 0, 0) FANOUT_792 (N7998, {N7998_0, N7998_1});
fanout_n #(2, 0, 0) FANOUT_793 (N8001, {N8001_0, N8001_1});
fanout_n #(2, 0, 0) FANOUT_794 (N8004, {N8004_0, N8004_1});
fanout_n #(2, 0, 0) FANOUT_795 (N8013, {N8013_0, N8013_1});
fanout_n #(2, 0, 0) FANOUT_796 (N8017, {N8017_0, N8017_1});
fanout_n #(2, 0, 0) FANOUT_797 (N8045, {N8045_0, N8045_1});
fanout_n #(2, 0, 0) FANOUT_798 (N8048, {N8048_0, N8048_1});
fanout_n #(2, 0, 0) FANOUT_799 (N8061, {N8061_0, N8061_1});
fanout_n #(2, 0, 0) FANOUT_800 (N8064, {N8064_0, N8064_1});
fanout_n #(2, 0, 0) FANOUT_801 (N8079, {N8079_0, N8079_1});
fanout_n #(2, 0, 0) FANOUT_802 (N8082, {N8082_0, N8082_1});
fanout_n #(2, 0, 0) FANOUT_803 (N8093, {N8093_0, N8093_1});
fanout_n #(2, 0, 0) FANOUT_804 (N8096, {N8096_0, N8096_1});
fanout_n #(2, 0, 0) FANOUT_805 (N8099, {N8099_0, N8099_1});
fanout_n #(2, 0, 0) FANOUT_806 (N8102, {N8102_0, N8102_1});


bufg #(0, 0) BUF_1 (N709, N141_0);
bufg #(0, 0) BUF_2 (N816, N293_0);
and_n #(2, 0, 0) AND_1 (N1042, {N135, N631});
notg #(0, 0) NOT_1 (N1043, N591);
bufg #(0, 0) BUF_3 (N1066, N592_0);
notg #(0, 0) NOT_2 (N1067, N595);
notg #(0, 0) NOT_3 (N1080, N596);
notg #(0, 0) NOT_4 (N1092, N597);
notg #(0, 0) NOT_5 (N1104, N598);
notg #(0, 0) NOT_6 (N1137, N545_0);
notg #(0, 0) NOT_7 (N1138, N348_0);
notg #(0, 0) NOT_8 (N1139, N366_0);
and_n #(2, 0, 0) AND_2 (N1140, {N552_0, N562_0});
notg #(0, 0) NOT_9 (N1141, N549_0);
notg #(0, 0) NOT_10 (N1142, N545_1);
notg #(0, 0) NOT_11 (N1143, N545_2);
notg #(0, 0) NOT_12 (N1144, N338_0);
notg #(0, 0) NOT_13 (N1145, N358_0);
nand_n #(2, 0, 0) NAND_1 (N1146, {N373, N1_0});
and_n #(2, 0, 0) AND_3 (N1147, {N141_1, N145});
notg #(0, 0) NOT_14 (N1148, N592_1);
notg #(0, 0) NOT_15 (N1149, N1042);
and_n #(2, 0, 0) AND_4 (N1150, {N1043, N27_0});
and_n #(2, 0, 0) AND_5 (N1151, {N386_0, N556_0});
notg #(0, 0) NOT_16 (N1152, N245_0);
notg #(0, 0) NOT_17 (N1153, N552_1);
notg #(0, 0) NOT_18 (N1154, N562_1);
notg #(0, 0) NOT_19 (N1155, N559_0);
and_n #(4, 0, 0) AND_6 (N1156, {N386_1, N559_1, N556_1, N552_2});
notg #(0, 0) NOT_20 (N1157, N566_0);
bufg #(0, 0) BUF_4 (N1161, N571_0);
bufg #(0, 0) BUF_5 (N1173, N574_0);
bufg #(0, 0) BUF_6 (N1185, N571_1);
bufg #(0, 0) BUF_7 (N1197, N574_1);
bufg #(0, 0) BUF_8 (N1209, N137_0);
bufg #(0, 0) BUF_9 (N1213, N137_1);
bufg #(0, 0) BUF_10 (N1216, N141_2);
notg #(0, 0) NOT_21 (N1219, N583_0);
bufg #(0, 0) BUF_11 (N1223, N577_0);
bufg #(0, 0) BUF_12 (N1235, N580_0);
bufg #(0, 0) BUF_13 (N1247, N577_1);
bufg #(0, 0) BUF_14 (N1259, N580_1);
bufg #(0, 0) BUF_15 (N1271, N254_0);
bufg #(0, 0) BUF_16 (N1280, N251_0);
bufg #(0, 0) BUF_17 (N1292, N251_1);
bufg #(0, 0) BUF_18 (N1303, N248_0);
bufg #(0, 0) BUF_19 (N1315, N248_1);
bufg #(0, 0) BUF_20 (N1327, N610_0);
bufg #(0, 0) BUF_21 (N1339, N607_0);
bufg #(0, 0) BUF_22 (N1351, N613_0);
bufg #(0, 0) BUF_23 (N1363, N616_0);
bufg #(0, 0) BUF_24 (N1375, N210_0);
bufg #(0, 0) BUF_25 (N1378, N210_1);
bufg #(0, 0) BUF_26 (N1381, N218_0);
bufg #(0, 0) BUF_27 (N1384, N218_1);
bufg #(0, 0) BUF_28 (N1387, N226_0);
bufg #(0, 0) BUF_29 (N1390, N226_1);
bufg #(0, 0) BUF_30 (N1393, N234_0);
bufg #(0, 0) BUF_31 (N1396, N234_1);
bufg #(0, 0) BUF_32 (N1415, N257_0);
bufg #(0, 0) BUF_33 (N1418, N257_1);
bufg #(0, 0) BUF_34 (N1421, N265_0);
bufg #(0, 0) BUF_35 (N1424, N265_1);
bufg #(0, 0) BUF_36 (N1427, N273_0);
bufg #(0, 0) BUF_37 (N1430, N273_1);
bufg #(0, 0) BUF_38 (N1433, N281_0);
bufg #(0, 0) BUF_39 (N1436, N281_1);
bufg #(0, 0) BUF_40 (N1455, N335_0);
bufg #(0, 0) BUF_41 (N1462, N335_1);
bufg #(0, 0) BUF_42 (N1469, N206_0);
and_n #(2, 0, 0) AND_7 (N1475, {N27_1, N31_0});
bufg #(0, 0) BUF_43 (N1479, N1_1);
bufg #(0, 0) BUF_44 (N1482, N588_0);
bufg #(0, 0) BUF_45 (N1492, N293_1);
bufg #(0, 0) BUF_46 (N1495, N302_0);
bufg #(0, 0) BUF_47 (N1498, N308_0);
bufg #(0, 0) BUF_48 (N1501, N308_1);
bufg #(0, 0) BUF_49 (N1504, N316_0);
bufg #(0, 0) BUF_50 (N1507, N316_1);
bufg #(0, 0) BUF_51 (N1510, N324_0);
bufg #(0, 0) BUF_52 (N1513, N324_1);
bufg #(0, 0) BUF_53 (N1516, N341_0);
bufg #(0, 0) BUF_54 (N1519, N341_1);
bufg #(0, 0) BUF_55 (N1522, N351_0);
bufg #(0, 0) BUF_56 (N1525, N351_1);
bufg #(0, 0) BUF_57 (N1542, N257_2);
bufg #(0, 0) BUF_58 (N1545, N257_3);
bufg #(0, 0) BUF_59 (N1548, N265_2);
bufg #(0, 0) BUF_60 (N1551, N265_3);
bufg #(0, 0) BUF_61 (N1554, N273_2);
bufg #(0, 0) BUF_62 (N1557, N273_3);
bufg #(0, 0) BUF_63 (N1560, N281_2);
bufg #(0, 0) BUF_64 (N1563, N281_3);
bufg #(0, 0) BUF_65 (N1566, N332_0);
bufg #(0, 0) BUF_66 (N1573, N332_1);
bufg #(0, 0) BUF_67 (N1580, N549_1);
and_n #(2, 0, 0) AND_8 (N1583, {N31_1, N27_2});
notg #(0, 0) NOT_22 (N1588, N588_1);
bufg #(0, 0) BUF_68 (N1594, N324_2);
bufg #(0, 0) BUF_69 (N1597, N324_3);
bufg #(0, 0) BUF_70 (N1600, N341_2);
bufg #(0, 0) BUF_71 (N1603, N341_3);
bufg #(0, 0) BUF_72 (N1606, N351_2);
bufg #(0, 0) BUF_73 (N1609, N351_3);
bufg #(0, 0) BUF_74 (N1612, N293_2);
bufg #(0, 0) BUF_75 (N1615, N302_1);
bufg #(0, 0) BUF_76 (N1618, N308_2);
bufg #(0, 0) BUF_77 (N1621, N308_3);
bufg #(0, 0) BUF_78 (N1624, N316_2);
bufg #(0, 0) BUF_79 (N1627, N316_3);
bufg #(0, 0) BUF_80 (N1630, N361_0);
bufg #(0, 0) BUF_81 (N1633, N361_1);
bufg #(0, 0) BUF_82 (N1636, N210_2);
bufg #(0, 0) BUF_83 (N1639, N210_3);
bufg #(0, 0) BUF_84 (N1642, N218_2);
bufg #(0, 0) BUF_85 (N1645, N218_3);
bufg #(0, 0) BUF_86 (N1648, N226_2);
bufg #(0, 0) BUF_87 (N1651, N226_3);
bufg #(0, 0) BUF_88 (N1654, N234_2);
bufg #(0, 0) BUF_89 (N1657, N234_3);
notg #(0, 0) NOT_23 (N1660, N324_4);
bufg #(0, 0) BUF_90 (N1663, N242_0);
bufg #(0, 0) BUF_91 (N1675, N242_1);
bufg #(0, 0) BUF_92 (N1685, N254_1);
bufg #(0, 0) BUF_93 (N1697, N610_1);
bufg #(0, 0) BUF_94 (N1709, N607_1);
bufg #(0, 0) BUF_95 (N1721, N625_0);
bufg #(0, 0) BUF_96 (N1727, N619_0);
bufg #(0, 0) BUF_97 (N1731, N613_1);
bufg #(0, 0) BUF_98 (N1743, N616_1);
notg #(0, 0) NOT_24 (N1755, N599_0);
notg #(0, 0) NOT_25 (N1758, N603_0);
bufg #(0, 0) BUF_99 (N1761, N619_1);
bufg #(0, 0) BUF_100 (N1769, N625_1);
bufg #(0, 0) BUF_101 (N1777, N619_2);
bufg #(0, 0) BUF_102 (N1785, N625_2);
bufg #(0, 0) BUF_103 (N1793, N619_3);
bufg #(0, 0) BUF_104 (N1800, N625_3);
bufg #(0, 0) BUF_105 (N1807, N619_4);
bufg #(0, 0) BUF_106 (N1814, N625_4);
bufg #(0, 0) BUF_107 (N1821, N299_0);
bufg #(0, 0) BUF_108 (N1824, N446_0);
bufg #(0, 0) BUF_109 (N1827, N457_0);
bufg #(0, 0) BUF_110 (N1830, N468_0);
bufg #(0, 0) BUF_111 (N1833, N422_0);
bufg #(0, 0) BUF_112 (N1836, N435_0);
bufg #(0, 0) BUF_113 (N1839, N389_0);
bufg #(0, 0) BUF_114 (N1842, N400_0);
bufg #(0, 0) BUF_115 (N1845, N411_0);
bufg #(0, 0) BUF_116 (N1848, N374_0);
bufg #(0, 0) BUF_117 (N1851, N4_0);
bufg #(0, 0) BUF_118 (N1854, N446_1);
bufg #(0, 0) BUF_119 (N1857, N457_1);
bufg #(0, 0) BUF_120 (N1860, N468_1);
bufg #(0, 0) BUF_121 (N1863, N435_1);
bufg #(0, 0) BUF_122 (N1866, N389_1);
bufg #(0, 0) BUF_123 (N1869, N400_1);
bufg #(0, 0) BUF_124 (N1872, N411_1);
bufg #(0, 0) BUF_125 (N1875, N422_1);
bufg #(0, 0) BUF_126 (N1878, N374_1);
bufg #(0, 0) BUF_127 (N1881, N479_0);
bufg #(0, 0) BUF_128 (N1884, N490_0);
bufg #(0, 0) BUF_129 (N1887, N503_0);
bufg #(0, 0) BUF_130 (N1890, N514_0);
bufg #(0, 0) BUF_131 (N1893, N523_0);
bufg #(0, 0) BUF_132 (N1896, N534_0);
bufg #(0, 0) BUF_133 (N1899, N54_0);
bufg #(0, 0) BUF_134 (N1902, N479_1);
bufg #(0, 0) BUF_135 (N1905, N503_1);
bufg #(0, 0) BUF_136 (N1908, N514_1);
bufg #(0, 0) BUF_137 (N1911, N523_1);
bufg #(0, 0) BUF_138 (N1914, N534_1);
bufg #(0, 0) BUF_139 (N1917, N490_1);
bufg #(0, 0) BUF_140 (N1920, N361_2);
bufg #(0, 0) BUF_141 (N1923, N369_0);
bufg #(0, 0) BUF_142 (N1926, N341_4);
bufg #(0, 0) BUF_143 (N1929, N351_4);
bufg #(0, 0) BUF_144 (N1932, N308_4);
bufg #(0, 0) BUF_145 (N1935, N316_4);
bufg #(0, 0) BUF_146 (N1938, N293_3);
bufg #(0, 0) BUF_147 (N1941, N302_2);
bufg #(0, 0) BUF_148 (N1944, N281_4);
bufg #(0, 0) BUF_149 (N1947, N289_0);
bufg #(0, 0) BUF_150 (N1950, N265_4);
bufg #(0, 0) BUF_151 (N1953, N273_4);
bufg #(0, 0) BUF_152 (N1956, N234_4);
bufg #(0, 0) BUF_153 (N1959, N257_4);
bufg #(0, 0) BUF_154 (N1962, N218_4);
bufg #(0, 0) BUF_155 (N1965, N226_4);
bufg #(0, 0) BUF_156 (N1968, N210_4);
notg #(0, 0) NOT_26 (N1972, N1146);
and_n #(2, 0, 0) AND_9 (N2054, {N136, N1148});
notg #(0, 0) NOT_27 (N2060, N1150);
notg #(0, 0) NOT_28 (N2061, N1151);
bufg #(0, 0) BUF_157 (N2139, N1209_0);
bufg #(0, 0) BUF_158 (N2142, N1216_0);
bufg #(0, 0) BUF_159 (N2309, N1479_0);
and_n #(2, 0, 0) AND_10 (N2349, {N1104_0, N514_2});
or_n #(2, 0, 0) OR_1 (N2350, {N1067_0, N514_3});
bufg #(0, 0) BUF_160 (N2387, N1580_0);
bufg #(0, 0) BUF_161 (N2527, N1821_0);
notg #(0, 0) NOT_29 (N2584, N1580_1);
and_n #(3, 0, 0) AND_11 (N2585, {N170_0, N1161_0, N1173_0});
and_n #(3, 0, 0) AND_12 (N2586, {N173_0, N1161_1, N1173_1});
and_n #(3, 0, 0) AND_13 (N2587, {N167_0, N1161_2, N1173_2});
and_n #(3, 0, 0) AND_14 (N2588, {N164_0, N1161_3, N1173_3});
and_n #(3, 0, 0) AND_15 (N2589, {N161_0, N1161_4, N1173_4});
nand_n #(2, 0, 0) NAND_2 (N2590, {N1475_0, N140});
and_n #(3, 0, 0) AND_16 (N2591, {N185_0, N1185_0, N1197_0});
and_n #(3, 0, 0) AND_17 (N2592, {N158_0, N1185_1, N1197_1});
and_n #(3, 0, 0) AND_18 (N2593, {N152_0, N1185_2, N1197_2});
and_n #(3, 0, 0) AND_19 (N2594, {N146_0, N1185_3, N1197_3});
and_n #(3, 0, 0) AND_20 (N2595, {N170_1, N1223_0, N1235_0});
and_n #(3, 0, 0) AND_21 (N2596, {N173_1, N1223_1, N1235_1});
and_n #(3, 0, 0) AND_22 (N2597, {N167_1, N1223_2, N1235_2});
and_n #(3, 0, 0) AND_23 (N2598, {N164_1, N1223_3, N1235_3});
and_n #(3, 0, 0) AND_24 (N2599, {N161_1, N1223_4, N1235_4});
and_n #(3, 0, 0) AND_25 (N2600, {N185_1, N1247_0, N1259_0});
and_n #(3, 0, 0) AND_26 (N2601, {N158_1, N1247_1, N1259_1});
and_n #(3, 0, 0) AND_27 (N2602, {N152_1, N1247_2, N1259_2});
and_n #(3, 0, 0) AND_28 (N2603, {N146_1, N1247_3, N1259_3});
and_n #(3, 0, 0) AND_29 (N2604, {N106_0, N1731_0, N1743_0});
and_n #(3, 0, 0) AND_30 (N2605, {N61_0, N1327_0, N1339_0});
and_n #(3, 0, 0) AND_31 (N2606, {N106_1, N1697_0, N1709_0});
and_n #(3, 0, 0) AND_32 (N2607, {N49_0, N1697_1, N1709_1});
and_n #(3, 0, 0) AND_33 (N2608, {N103_0, N1697_2, N1709_2});
and_n #(3, 0, 0) AND_34 (N2609, {N40_0, N1697_3, N1709_3});
and_n #(3, 0, 0) AND_35 (N2610, {N37_0, N1697_4, N1709_4});
and_n #(3, 0, 0) AND_36 (N2611, {N20_0, N1327_1, N1339_1});
and_n #(3, 0, 0) AND_37 (N2612, {N17_0, N1327_2, N1339_2});
and_n #(3, 0, 0) AND_38 (N2613, {N70_0, N1327_3, N1339_3});
and_n #(3, 0, 0) AND_39 (N2614, {N64_0, N1327_4, N1339_4});
and_n #(3, 0, 0) AND_40 (N2615, {N49_1, N1731_1, N1743_1});
and_n #(3, 0, 0) AND_41 (N2616, {N103_1, N1731_2, N1743_2});
and_n #(3, 0, 0) AND_42 (N2617, {N40_1, N1731_3, N1743_3});
and_n #(3, 0, 0) AND_43 (N2618, {N37_1, N1731_4, N1743_4});
and_n #(3, 0, 0) AND_44 (N2619, {N20_1, N1351_0, N1363_0});
and_n #(3, 0, 0) AND_45 (N2620, {N17_1, N1351_1, N1363_1});
and_n #(3, 0, 0) AND_46 (N2621, {N70_1, N1351_2, N1363_2});
and_n #(3, 0, 0) AND_47 (N2622, {N64_1, N1351_3, N1363_3});
notg #(0, 0) NOT_30 (N2623, N1475_1);
and_n #(3, 0, 0) AND_48 (N2624, {N123_0, N1758_0, N599_1});
and_n #(2, 0, 0) AND_49 (N2625, {N1777_0, N1785_0});
and_n #(3, 0, 0) AND_50 (N2626, {N61_1, N1351_4, N1363_4});
and_n #(2, 0, 0) AND_51 (N2627, {N1761_0, N1769_0});
notg #(0, 0) NOT_31 (N2628, N1824_0);
notg #(0, 0) NOT_32 (N2629, N1827_0);
notg #(0, 0) NOT_33 (N2630, N1830_0);
notg #(0, 0) NOT_34 (N2631, N1833_0);
notg #(0, 0) NOT_35 (N2632, N1836_0);
notg #(0, 0) NOT_36 (N2633, N1839_0);
notg #(0, 0) NOT_37 (N2634, N1842_0);
notg #(0, 0) NOT_38 (N2635, N1845_0);
notg #(0, 0) NOT_39 (N2636, N1848_0);
notg #(0, 0) NOT_40 (N2637, N1851_0);
notg #(0, 0) NOT_41 (N2638, N1854_0);
notg #(0, 0) NOT_42 (N2639, N1857_0);
notg #(0, 0) NOT_43 (N2640, N1860_0);
notg #(0, 0) NOT_44 (N2641, N1863_0);
notg #(0, 0) NOT_45 (N2642, N1866_0);
notg #(0, 0) NOT_46 (N2643, N1869_0);
notg #(0, 0) NOT_47 (N2644, N1872_0);
notg #(0, 0) NOT_48 (N2645, N1875_0);
notg #(0, 0) NOT_49 (N2646, N1878_0);
bufg #(0, 0) BUF_162 (N2647, N1209_1);
notg #(0, 0) NOT_50 (N2653, N1161_5);
notg #(0, 0) NOT_51 (N2664, N1173_5);
bufg #(0, 0) BUF_163 (N2675, N1209_2);
notg #(0, 0) NOT_52 (N2681, N1185_4);
notg #(0, 0) NOT_53 (N2692, N1197_4);
and_n #(3, 0, 0) AND_52 (N2703, {N179_0, N1185_5, N1197_5});
bufg #(0, 0) BUF_164 (N2704, N1479_1);
notg #(0, 0) NOT_54 (N2709, N1881_0);
notg #(0, 0) NOT_55 (N2710, N1884_0);
notg #(0, 0) NOT_56 (N2711, N1887_0);
notg #(0, 0) NOT_57 (N2712, N1890_0);
notg #(0, 0) NOT_58 (N2713, N1893_0);
notg #(0, 0) NOT_59 (N2714, N1896_0);
notg #(0, 0) NOT_60 (N2715, N1899_0);
notg #(0, 0) NOT_61 (N2716, N1902_0);
notg #(0, 0) NOT_62 (N2717, N1905_0);
notg #(0, 0) NOT_63 (N2718, N1908_0);
notg #(0, 0) NOT_64 (N2719, N1911_0);
notg #(0, 0) NOT_65 (N2720, N1914_0);
notg #(0, 0) NOT_66 (N2721, N1917_0);
bufg #(0, 0) BUF_165 (N2722, N1213_0);
notg #(0, 0) NOT_67 (N2728, N1223_5);
notg #(0, 0) NOT_68 (N2739, N1235_5);
bufg #(0, 0) BUF_166 (N2750, N1213_1);
notg #(0, 0) NOT_69 (N2756, N1247_4);
notg #(0, 0) NOT_70 (N2767, N1259_4);
and_n #(3, 0, 0) AND_53 (N2778, {N179_1, N1247_5, N1259_5});
notg #(0, 0) NOT_71 (N2779, N1327_5);
notg #(0, 0) NOT_72 (N2790, N1339_5);
notg #(0, 0) NOT_73 (N2801, N1351_5);
notg #(0, 0) NOT_74 (N2812, N1363_5);
notg #(0, 0) NOT_75 (N2823, N1375_0);
notg #(0, 0) NOT_76 (N2824, N1378_0);
notg #(0, 0) NOT_77 (N2825, N1381_0);
notg #(0, 0) NOT_78 (N2826, N1384_0);
notg #(0, 0) NOT_79 (N2827, N1387_0);
notg #(0, 0) NOT_80 (N2828, N1390_0);
notg #(0, 0) NOT_81 (N2829, N1393_0);
notg #(0, 0) NOT_82 (N2830, N1396_0);
and_n #(3, 0, 0) AND_54 (N2831, {N1104_1, N457_2, N1378_1});
and_n #(3, 0, 0) AND_55 (N2832, {N1104_2, N468_2, N1384_1});
and_n #(3, 0, 0) AND_56 (N2833, {N1104_3, N422_2, N1390_1});
and_n #(3, 0, 0) AND_57 (N2834, {N1104_4, N435_2, N1396_1});
and_n #(2, 0, 0) AND_58 (N2835, {N1067_1, N1375_1});
and_n #(2, 0, 0) AND_59 (N2836, {N1067_2, N1381_1});
and_n #(2, 0, 0) AND_60 (N2837, {N1067_3, N1387_1});
and_n #(2, 0, 0) AND_61 (N2838, {N1067_4, N1393_1});
notg #(0, 0) NOT_83 (N2839, N1415_0);
notg #(0, 0) NOT_84 (N2840, N1418_0);
notg #(0, 0) NOT_85 (N2841, N1421_0);
notg #(0, 0) NOT_86 (N2842, N1424_0);
notg #(0, 0) NOT_87 (N2843, N1427_0);
notg #(0, 0) NOT_88 (N2844, N1430_0);
notg #(0, 0) NOT_89 (N2845, N1433_0);
notg #(0, 0) NOT_90 (N2846, N1436_0);
and_n #(3, 0, 0) AND_62 (N2847, {N1104_5, N389_2, N1418_1});
and_n #(3, 0, 0) AND_63 (N2848, {N1104_6, N400_2, N1424_1});
and_n #(3, 0, 0) AND_64 (N2849, {N1104_7, N411_2, N1430_1});
and_n #(3, 0, 0) AND_65 (N2850, {N1104_8, N374_2, N1436_1});
and_n #(2, 0, 0) AND_66 (N2851, {N1067_5, N1415_1});
and_n #(2, 0, 0) AND_67 (N2852, {N1067_6, N1421_1});
and_n #(2, 0, 0) AND_68 (N2853, {N1067_7, N1427_1});
and_n #(2, 0, 0) AND_69 (N2854, {N1067_8, N1433_1});
notg #(0, 0) NOT_91 (N2855, N1455_0);
notg #(0, 0) NOT_92 (N2861, N1462_0);
and_n #(2, 0, 0) AND_70 (N2867, {N292, N1455_1});
and_n #(2, 0, 0) AND_71 (N2868, {N288, N1455_2});
and_n #(2, 0, 0) AND_72 (N2869, {N280, N1455_3});
and_n #(2, 0, 0) AND_73 (N2870, {N272, N1455_4});
and_n #(2, 0, 0) AND_74 (N2871, {N264, N1455_5});
and_n #(2, 0, 0) AND_75 (N2872, {N241, N1462_1});
and_n #(2, 0, 0) AND_76 (N2873, {N233, N1462_2});
and_n #(2, 0, 0) AND_77 (N2874, {N225, N1462_3});
and_n #(2, 0, 0) AND_78 (N2875, {N217, N1462_4});
and_n #(2, 0, 0) AND_79 (N2876, {N209, N1462_5});
bufg #(0, 0) BUF_167 (N2877, N1216_1);
notg #(0, 0) NOT_93 (N2882, N1482_0);
notg #(0, 0) NOT_94 (N2891, N1475_2);
notg #(0, 0) NOT_95 (N2901, N1492_0);
notg #(0, 0) NOT_96 (N2902, N1495_0);
notg #(0, 0) NOT_97 (N2903, N1498_0);
notg #(0, 0) NOT_98 (N2904, N1501_0);
notg #(0, 0) NOT_99 (N2905, N1504_0);
notg #(0, 0) NOT_100 (N2906, N1507_0);
and_n #(2, 0, 0) AND_80 (N2907, {N1303_0, N1495_1});
and_n #(3, 0, 0) AND_81 (N2908, {N1303_1, N479_2, N1501_1});
and_n #(3, 0, 0) AND_82 (N2909, {N1303_2, N490_2, N1507_1});
and_n #(2, 0, 0) AND_83 (N2910, {N1663_0, N1492_1});
and_n #(2, 0, 0) AND_84 (N2911, {N1663_1, N1498_1});
and_n #(2, 0, 0) AND_85 (N2912, {N1663_2, N1504_1});
notg #(0, 0) NOT_101 (N2913, N1510_0);
notg #(0, 0) NOT_102 (N2914, N1513_0);
notg #(0, 0) NOT_103 (N2915, N1516_0);
notg #(0, 0) NOT_104 (N2916, N1519_0);
notg #(0, 0) NOT_105 (N2917, N1522_0);
notg #(0, 0) NOT_106 (N2918, N1525_0);
and_n #(3, 0, 0) AND_86 (N2919, {N1104_9, N503_2, N1513_1});
notg #(0, 0) NOT_107 (N2920, N2349);
and_n #(3, 0, 0) AND_87 (N2921, {N1104_10, N523_2, N1519_1});
and_n #(3, 0, 0) AND_88 (N2922, {N1104_11, N534_2, N1525_1});
and_n #(2, 0, 0) AND_89 (N2923, {N1067_9, N1510_1});
and_n #(2, 0, 0) AND_90 (N2924, {N1067_10, N1516_1});
and_n #(2, 0, 0) AND_91 (N2925, {N1067_11, N1522_1});
notg #(0, 0) NOT_108 (N2926, N1542_0);
notg #(0, 0) NOT_109 (N2927, N1545_0);
notg #(0, 0) NOT_110 (N2928, N1548_0);
notg #(0, 0) NOT_111 (N2929, N1551_0);
notg #(0, 0) NOT_112 (N2930, N1554_0);
notg #(0, 0) NOT_113 (N2931, N1557_0);
notg #(0, 0) NOT_114 (N2932, N1560_0);
notg #(0, 0) NOT_115 (N2933, N1563_0);
and_n #(3, 0, 0) AND_92 (N2934, {N1303_3, N389_3, N1545_1});
and_n #(3, 0, 0) AND_93 (N2935, {N1303_4, N400_3, N1551_1});
and_n #(3, 0, 0) AND_94 (N2936, {N1303_5, N411_3, N1557_1});
and_n #(3, 0, 0) AND_95 (N2937, {N1303_6, N374_3, N1563_1});
and_n #(2, 0, 0) AND_96 (N2938, {N1663_3, N1542_1});
and_n #(2, 0, 0) AND_97 (N2939, {N1663_4, N1548_1});
and_n #(2, 0, 0) AND_98 (N2940, {N1663_5, N1554_1});
and_n #(2, 0, 0) AND_99 (N2941, {N1663_6, N1560_1});
notg #(0, 0) NOT_116 (N2942, N1566_0);
notg #(0, 0) NOT_117 (N2948, N1573_0);
and_n #(2, 0, 0) AND_100 (N2954, {N372, N1566_1});
and_n #(2, 0, 0) AND_101 (N2955, {N366_1, N1566_2});
and_n #(2, 0, 0) AND_102 (N2956, {N358_1, N1566_3});
and_n #(2, 0, 0) AND_103 (N2957, {N348_1, N1566_4});
and_n #(2, 0, 0) AND_104 (N2958, {N338_1, N1566_5});
and_n #(2, 0, 0) AND_105 (N2959, {N331, N1573_1});
and_n #(2, 0, 0) AND_106 (N2960, {N323, N1573_2});
and_n #(2, 0, 0) AND_107 (N2961, {N315, N1573_3});
and_n #(2, 0, 0) AND_108 (N2962, {N307, N1573_4});
and_n #(2, 0, 0) AND_109 (N2963, {N299_1, N1573_5});
notg #(0, 0) NOT_118 (N2964, N1588_0);
and_n #(2, 0, 0) AND_110 (N2969, {N83_0, N1588_1});
and_n #(2, 0, 0) AND_111 (N2970, {N86, N1588_2});
and_n #(2, 0, 0) AND_112 (N2971, {N88_0, N1588_3});
and_n #(2, 0, 0) AND_113 (N2972, {N88_1, N1588_4});
notg #(0, 0) NOT_119 (N2973, N1594_0);
notg #(0, 0) NOT_120 (N2974, N1597_0);
notg #(0, 0) NOT_121 (N2975, N1600_0);
notg #(0, 0) NOT_122 (N2976, N1603_0);
notg #(0, 0) NOT_123 (N2977, N1606_0);
notg #(0, 0) NOT_124 (N2978, N1609_0);
and_n #(3, 0, 0) AND_114 (N2979, {N1315_0, N503_3, N1597_1});
and_n #(2, 0, 0) AND_115 (N2980, {N1315_1, N514_4});
and_n #(3, 0, 0) AND_116 (N2981, {N1315_2, N523_3, N1603_1});
and_n #(3, 0, 0) AND_117 (N2982, {N1315_3, N534_3, N1609_1});
and_n #(2, 0, 0) AND_118 (N2983, {N1675_0, N1594_1});
or_n #(2, 0, 0) OR_2 (N2984, {N1675_1, N514_5});
and_n #(2, 0, 0) AND_119 (N2985, {N1675_2, N1600_1});
and_n #(2, 0, 0) AND_120 (N2986, {N1675_3, N1606_1});
notg #(0, 0) NOT_125 (N2987, N1612_0);
notg #(0, 0) NOT_126 (N2988, N1615_0);
notg #(0, 0) NOT_127 (N2989, N1618_0);
notg #(0, 0) NOT_128 (N2990, N1621_0);
notg #(0, 0) NOT_129 (N2991, N1624_0);
notg #(0, 0) NOT_130 (N2992, N1627_0);
and_n #(2, 0, 0) AND_121 (N2993, {N1315_4, N1615_1});
and_n #(3, 0, 0) AND_122 (N2994, {N1315_5, N479_3, N1621_1});
and_n #(3, 0, 0) AND_123 (N2995, {N1315_6, N490_3, N1627_1});
and_n #(2, 0, 0) AND_124 (N2996, {N1675_4, N1612_1});
and_n #(2, 0, 0) AND_125 (N2997, {N1675_5, N1618_1});
and_n #(2, 0, 0) AND_126 (N2998, {N1675_6, N1624_1});
notg #(0, 0) NOT_131 (N2999, N1630_0);
bufg #(0, 0) BUF_168 (N3000, N1469_0);
bufg #(0, 0) BUF_169 (N3003, N1469_1);
notg #(0, 0) NOT_132 (N3006, N1633_0);
bufg #(0, 0) BUF_170 (N3007, N1469_2);
bufg #(0, 0) BUF_171 (N3010, N1469_3);
and_n #(2, 0, 0) AND_127 (N3013, {N1315_7, N1630_1});
and_n #(2, 0, 0) AND_128 (N3014, {N1315_8, N1633_1});
notg #(0, 0) NOT_133 (N3015, N1636_0);
notg #(0, 0) NOT_134 (N3016, N1639_0);
notg #(0, 0) NOT_135 (N3017, N1642_0);
notg #(0, 0) NOT_136 (N3018, N1645_0);
notg #(0, 0) NOT_137 (N3019, N1648_0);
notg #(0, 0) NOT_138 (N3020, N1651_0);
notg #(0, 0) NOT_139 (N3021, N1654_0);
notg #(0, 0) NOT_140 (N3022, N1657_0);
and_n #(3, 0, 0) AND_129 (N3023, {N1303_7, N457_3, N1639_1});
and_n #(3, 0, 0) AND_130 (N3024, {N1303_8, N468_3, N1645_1});
and_n #(3, 0, 0) AND_131 (N3025, {N1303_9, N422_3, N1651_1});
and_n #(3, 0, 0) AND_132 (N3026, {N1303_10, N435_3, N1657_1});
and_n #(2, 0, 0) AND_133 (N3027, {N1663_7, N1636_1});
and_n #(2, 0, 0) AND_134 (N3028, {N1663_8, N1642_1});
and_n #(2, 0, 0) AND_135 (N3029, {N1663_9, N1648_1});
and_n #(2, 0, 0) AND_136 (N3030, {N1663_10, N1654_1});
notg #(0, 0) NOT_141 (N3031, N1920_0);
notg #(0, 0) NOT_142 (N3032, N1923_0);
notg #(0, 0) NOT_143 (N3033, N1926_0);
notg #(0, 0) NOT_144 (N3034, N1929_0);
bufg #(0, 0) BUF_172 (N3035, N1660_0);
bufg #(0, 0) BUF_173 (N3038, N1660_1);
notg #(0, 0) NOT_145 (N3041, N1697_5);
notg #(0, 0) NOT_146 (N3052, N1709_5);
notg #(0, 0) NOT_147 (N3063, N1721_0);
notg #(0, 0) NOT_148 (N3068, N1727_0);
and_n #(2, 0, 0) AND_137 (N3071, {N97_0, N1721_1});
and_n #(2, 0, 0) AND_138 (N3072, {N94_0, N1721_2});
and_n #(2, 0, 0) AND_139 (N3073, {N97_1, N1721_3});
and_n #(2, 0, 0) AND_140 (N3074, {N94_1, N1721_4});
notg #(0, 0) NOT_149 (N3075, N1731_5);
notg #(0, 0) NOT_150 (N3086, N1743_5);
notg #(0, 0) NOT_151 (N3097, N1761_1);
notg #(0, 0) NOT_152 (N3108, N1769_1);
notg #(0, 0) NOT_153 (N3119, N1777_1);
notg #(0, 0) NOT_154 (N3130, N1785_1);
notg #(0, 0) NOT_155 (N3141, N1944_0);
notg #(0, 0) NOT_156 (N3142, N1947_0);
notg #(0, 0) NOT_157 (N3143, N1950_0);
notg #(0, 0) NOT_158 (N3144, N1953_0);
notg #(0, 0) NOT_159 (N3145, N1956_0);
notg #(0, 0) NOT_160 (N3146, N1959_0);
notg #(0, 0) NOT_161 (N3147, N1793_0);
notg #(0, 0) NOT_162 (N3158, N1800_0);
notg #(0, 0) NOT_163 (N3169, N1807_0);
notg #(0, 0) NOT_164 (N3180, N1814_0);
bufg #(0, 0) BUF_174 (N3191, N1821_1);
notg #(0, 0) NOT_165 (N3194, N1932_0);
notg #(0, 0) NOT_166 (N3195, N1935_0);
notg #(0, 0) NOT_167 (N3196, N1938_0);
notg #(0, 0) NOT_168 (N3197, N1941_0);
notg #(0, 0) NOT_169 (N3198, N1962_0);
notg #(0, 0) NOT_170 (N3199, N1965_0);
bufg #(0, 0) BUF_175 (N3200, N1469_4);
notg #(0, 0) NOT_171 (N3203, N1968_0);
bufg #(0, 0) BUF_176 (N3357, N2704_0);
bufg #(0, 0) BUF_177 (N3358, N2704_1);
bufg #(0, 0) BUF_178 (N3359, N2704_2);
bufg #(0, 0) BUF_179 (N3360, N2704_3);
and_n #(3, 0, 0) AND_141 (N3401, {N457_4, N1092_0, N2824});
and_n #(3, 0, 0) AND_142 (N3402, {N468_4, N1092_1, N2826});
and_n #(3, 0, 0) AND_143 (N3403, {N422_4, N1092_2, N2828});
and_n #(3, 0, 0) AND_144 (N3404, {N435_4, N1092_3, N2830});
and_n #(2, 0, 0) AND_145 (N3405, {N1080_0, N2823});
and_n #(2, 0, 0) AND_146 (N3406, {N1080_1, N2825});
and_n #(2, 0, 0) AND_147 (N3407, {N1080_2, N2827});
and_n #(2, 0, 0) AND_148 (N3408, {N1080_3, N2829});
and_n #(3, 0, 0) AND_149 (N3409, {N389_4, N1092_4, N2840});
and_n #(3, 0, 0) AND_150 (N3410, {N400_4, N1092_5, N2842});
and_n #(3, 0, 0) AND_151 (N3411, {N411_4, N1092_6, N2844});
and_n #(3, 0, 0) AND_152 (N3412, {N374_4, N1092_7, N2846});
and_n #(2, 0, 0) AND_153 (N3413, {N1080_4, N2839});
and_n #(2, 0, 0) AND_154 (N3414, {N1080_5, N2841});
and_n #(2, 0, 0) AND_155 (N3415, {N1080_6, N2843});
and_n #(2, 0, 0) AND_156 (N3416, {N1080_7, N2845});
and_n #(2, 0, 0) AND_157 (N3444, {N1280_0, N2902});
and_n #(3, 0, 0) AND_158 (N3445, {N479_4, N1280_1, N2904});
and_n #(3, 0, 0) AND_159 (N3446, {N490_4, N1280_2, N2906});
and_n #(2, 0, 0) AND_160 (N3447, {N1685_0, N2901});
and_n #(2, 0, 0) AND_161 (N3448, {N1685_1, N2903});
and_n #(2, 0, 0) AND_162 (N3449, {N1685_2, N2905});
and_n #(3, 0, 0) AND_163 (N3450, {N503_4, N1092_8, N2914});
and_n #(3, 0, 0) AND_164 (N3451, {N523_4, N1092_9, N2916});
and_n #(3, 0, 0) AND_165 (N3452, {N534_4, N1092_10, N2918});
and_n #(2, 0, 0) AND_166 (N3453, {N1080_8, N2913});
and_n #(2, 0, 0) AND_167 (N3454, {N1080_9, N2915});
and_n #(2, 0, 0) AND_168 (N3455, {N1080_10, N2917});
and_n #(2, 0, 0) AND_169 (N3456, {N2920, N2350});
and_n #(3, 0, 0) AND_170 (N3459, {N389_5, N1280_3, N2927});
and_n #(3, 0, 0) AND_171 (N3460, {N400_5, N1280_4, N2929});
and_n #(3, 0, 0) AND_172 (N3461, {N411_5, N1280_5, N2931});
and_n #(3, 0, 0) AND_173 (N3462, {N374_5, N1280_6, N2933});
and_n #(2, 0, 0) AND_174 (N3463, {N1685_3, N2926});
and_n #(2, 0, 0) AND_175 (N3464, {N1685_4, N2928});
and_n #(2, 0, 0) AND_176 (N3465, {N1685_5, N2930});
and_n #(2, 0, 0) AND_177 (N3466, {N1685_6, N2932});
and_n #(3, 0, 0) AND_178 (N3481, {N503_5, N1292_0, N2974});
notg #(0, 0) NOT_172 (N3482, N2980);
and_n #(3, 0, 0) AND_179 (N3483, {N523_5, N1292_1, N2976});
and_n #(3, 0, 0) AND_180 (N3484, {N534_5, N1292_2, N2978});
and_n #(2, 0, 0) AND_181 (N3485, {N1271_0, N2973});
and_n #(2, 0, 0) AND_182 (N3486, {N1271_1, N2975});
and_n #(2, 0, 0) AND_183 (N3487, {N1271_2, N2977});
and_n #(2, 0, 0) AND_184 (N3488, {N1292_3, N2988});
and_n #(3, 0, 0) AND_185 (N3489, {N479_5, N1292_4, N2990});
and_n #(3, 0, 0) AND_186 (N3490, {N490_5, N1292_5, N2992});
and_n #(2, 0, 0) AND_187 (N3491, {N1271_3, N2987});
and_n #(2, 0, 0) AND_188 (N3492, {N1271_4, N2989});
and_n #(2, 0, 0) AND_189 (N3493, {N1271_5, N2991});
and_n #(2, 0, 0) AND_190 (N3502, {N1292_6, N2999});
and_n #(2, 0, 0) AND_191 (N3503, {N1292_7, N3006});
and_n #(3, 0, 0) AND_192 (N3504, {N457_5, N1280_7, N3016});
and_n #(3, 0, 0) AND_193 (N3505, {N468_5, N1280_8, N3018});
and_n #(3, 0, 0) AND_194 (N3506, {N422_5, N1280_9, N3020});
and_n #(3, 0, 0) AND_195 (N3507, {N435_5, N1280_10, N3022});
and_n #(2, 0, 0) AND_196 (N3508, {N1685_7, N3015});
and_n #(2, 0, 0) AND_197 (N3509, {N1685_8, N3017});
and_n #(2, 0, 0) AND_198 (N3510, {N1685_9, N3019});
and_n #(2, 0, 0) AND_199 (N3511, {N1685_10, N3021});
nand_n #(2, 0, 0) NAND_3 (N3512, {N1923_1, N3031});
nand_n #(2, 0, 0) NAND_4 (N3513, {N1920_1, N3032});
nand_n #(2, 0, 0) NAND_5 (N3514, {N1929_1, N3033});
nand_n #(2, 0, 0) NAND_6 (N3515, {N1926_1, N3034});
nand_n #(2, 0, 0) NAND_7 (N3558, {N1947_1, N3141});
nand_n #(2, 0, 0) NAND_8 (N3559, {N1944_1, N3142});
nand_n #(2, 0, 0) NAND_9 (N3560, {N1953_1, N3143});
nand_n #(2, 0, 0) NAND_10 (N3561, {N1950_1, N3144});
nand_n #(2, 0, 0) NAND_11 (N3562, {N1959_1, N3145});
nand_n #(2, 0, 0) NAND_12 (N3563, {N1956_1, N3146});
bufg #(0, 0) BUF_180 (N3604, N3191_0);
nand_n #(2, 0, 0) NAND_13 (N3605, {N1935_1, N3194});
nand_n #(2, 0, 0) NAND_14 (N3606, {N1932_1, N3195});
nand_n #(2, 0, 0) NAND_15 (N3607, {N1941_1, N3196});
nand_n #(2, 0, 0) NAND_16 (N3608, {N1938_1, N3197});
nand_n #(2, 0, 0) NAND_17 (N3609, {N1965_1, N3198});
nand_n #(2, 0, 0) NAND_18 (N3610, {N1962_1, N3199});
notg #(0, 0) NOT_173 (N3613, N3191_1);
and_n #(2, 0, 0) AND_200 (N3614, {N2882_0, N2891_0});
and_n #(2, 0, 0) AND_201 (N3615, {N1482_1, N2891_1});
and_n #(3, 0, 0) AND_202 (N3616, {N200_0, N2653_0, N1173_6});
and_n #(3, 0, 0) AND_203 (N3617, {N203_0, N2653_1, N1173_7});
and_n #(3, 0, 0) AND_204 (N3618, {N197_0, N2653_2, N1173_8});
and_n #(3, 0, 0) AND_205 (N3619, {N194_0, N2653_3, N1173_9});
and_n #(3, 0, 0) AND_206 (N3620, {N191_0, N2653_4, N1173_10});
and_n #(3, 0, 0) AND_207 (N3621, {N182_0, N2681_0, N1197_6});
and_n #(3, 0, 0) AND_208 (N3622, {N188_0, N2681_1, N1197_7});
and_n #(3, 0, 0) AND_209 (N3623, {N155_0, N2681_2, N1197_8});
and_n #(3, 0, 0) AND_210 (N3624, {N149_0, N2681_3, N1197_9});
and_n #(2, 0, 0) AND_211 (N3625, {N2882_1, N2891_2});
and_n #(2, 0, 0) AND_212 (N3626, {N1482_2, N2891_3});
and_n #(3, 0, 0) AND_213 (N3627, {N200_1, N2728_0, N1235_6});
and_n #(3, 0, 0) AND_214 (N3628, {N203_1, N2728_1, N1235_7});
and_n #(3, 0, 0) AND_215 (N3629, {N197_1, N2728_2, N1235_8});
and_n #(3, 0, 0) AND_216 (N3630, {N194_1, N2728_3, N1235_9});
and_n #(3, 0, 0) AND_217 (N3631, {N191_1, N2728_4, N1235_10});
and_n #(3, 0, 0) AND_218 (N3632, {N182_1, N2756_0, N1259_6});
and_n #(3, 0, 0) AND_219 (N3633, {N188_1, N2756_1, N1259_7});
and_n #(3, 0, 0) AND_220 (N3634, {N155_1, N2756_2, N1259_8});
and_n #(3, 0, 0) AND_221 (N3635, {N149_1, N2756_3, N1259_9});
and_n #(2, 0, 0) AND_222 (N3636, {N2882_2, N2891_4});
and_n #(2, 0, 0) AND_223 (N3637, {N1482_3, N2891_5});
and_n #(3, 0, 0) AND_224 (N3638, {N109_0, N3075_0, N1743_6});
and_n #(2, 0, 0) AND_225 (N3639, {N2882_3, N2891_6});
and_n #(2, 0, 0) AND_226 (N3640, {N1482_4, N2891_7});
and_n #(3, 0, 0) AND_227 (N3641, {N11_0, N2779_0, N1339_6});
and_n #(3, 0, 0) AND_228 (N3642, {N109_1, N3041_0, N1709_6});
and_n #(3, 0, 0) AND_229 (N3643, {N46_0, N3041_1, N1709_7});
and_n #(3, 0, 0) AND_230 (N3644, {N100_0, N3041_2, N1709_8});
and_n #(3, 0, 0) AND_231 (N3645, {N91_0, N3041_3, N1709_9});
and_n #(3, 0, 0) AND_232 (N3646, {N43_0, N3041_4, N1709_10});
and_n #(3, 0, 0) AND_233 (N3647, {N76_0, N2779_1, N1339_7});
and_n #(3, 0, 0) AND_234 (N3648, {N73_0, N2779_2, N1339_8});
and_n #(3, 0, 0) AND_235 (N3649, {N67_0, N2779_3, N1339_9});
and_n #(3, 0, 0) AND_236 (N3650, {N14_0, N2779_4, N1339_10});
and_n #(3, 0, 0) AND_237 (N3651, {N46_1, N3075_1, N1743_7});
and_n #(3, 0, 0) AND_238 (N3652, {N100_1, N3075_2, N1743_8});
and_n #(3, 0, 0) AND_239 (N3653, {N91_1, N3075_3, N1743_9});
and_n #(3, 0, 0) AND_240 (N3654, {N43_1, N3075_4, N1743_10});
and_n #(3, 0, 0) AND_241 (N3655, {N76_1, N2801_0, N1363_6});
and_n #(3, 0, 0) AND_242 (N3656, {N73_1, N2801_1, N1363_7});
and_n #(3, 0, 0) AND_243 (N3657, {N67_1, N2801_2, N1363_8});
and_n #(3, 0, 0) AND_244 (N3658, {N14_1, N2801_3, N1363_9});
and_n #(3, 0, 0) AND_245 (N3659, {N120, N3119_0, N1785_2});
and_n #(3, 0, 0) AND_246 (N3660, {N11_1, N2801_4, N1363_10});
and_n #(3, 0, 0) AND_247 (N3661, {N118, N3097_0, N1769_2});
and_n #(3, 0, 0) AND_248 (N3662, {N176_0, N2681_4, N1197_10});
and_n #(3, 0, 0) AND_249 (N3663, {N176_1, N2756_4, N1259_10});
or_n #(2, 0, 0) OR_3 (N3664, {N2831, N3401});
or_n #(2, 0, 0) OR_4 (N3665, {N2832, N3402});
or_n #(2, 0, 0) OR_5 (N3666, {N2833, N3403});
or_n #(2, 0, 0) OR_6 (N3667, {N2834, N3404});
or_n #(3, 0, 0) OR_7 (N3668, {N2835, N3405, N457_6});
or_n #(3, 0, 0) OR_8 (N3669, {N2836, N3406, N468_6});
or_n #(3, 0, 0) OR_9 (N3670, {N2837, N3407, N422_6});
or_n #(3, 0, 0) OR_10 (N3671, {N2838, N3408, N435_6});
or_n #(2, 0, 0) OR_11 (N3672, {N2847, N3409});
or_n #(2, 0, 0) OR_12 (N3673, {N2848, N3410});
or_n #(2, 0, 0) OR_13 (N3674, {N2849, N3411});
or_n #(2, 0, 0) OR_14 (N3675, {N2850, N3412});
or_n #(3, 0, 0) OR_15 (N3676, {N2851, N3413, N389_6});
or_n #(3, 0, 0) OR_16 (N3677, {N2852, N3414, N400_6});
or_n #(3, 0, 0) OR_17 (N3678, {N2853, N3415, N411_6});
or_n #(3, 0, 0) OR_18 (N3679, {N2854, N3416, N374_6});
and_n #(2, 0, 0) AND_250 (N3680, {N289_1, N2855_0});
and_n #(2, 0, 0) AND_251 (N3681, {N281_5, N2855_1});
and_n #(2, 0, 0) AND_252 (N3682, {N273_5, N2855_2});
and_n #(2, 0, 0) AND_253 (N3683, {N265_5, N2855_3});
and_n #(2, 0, 0) AND_254 (N3684, {N257_5, N2855_4});
and_n #(2, 0, 0) AND_255 (N3685, {N234_5, N2861_0});
and_n #(2, 0, 0) AND_256 (N3686, {N226_5, N2861_1});
and_n #(2, 0, 0) AND_257 (N3687, {N218_5, N2861_2});
and_n #(2, 0, 0) AND_258 (N3688, {N210_5, N2861_3});
and_n #(2, 0, 0) AND_259 (N3689, {N206_1, N2861_4});
notg #(0, 0) NOT_174 (N3691, N2891_8);
or_n #(2, 0, 0) OR_19 (N3700, {N2907, N3444});
or_n #(2, 0, 0) OR_20 (N3701, {N2908, N3445});
or_n #(2, 0, 0) OR_21 (N3702, {N2909, N3446});
or_n #(3, 0, 0) OR_22 (N3703, {N2911, N3448, N479_6});
or_n #(3, 0, 0) OR_23 (N3704, {N2912, N3449, N490_6});
or_n #(2, 0, 0) OR_24 (N3705, {N2910, N3447});
or_n #(2, 0, 0) OR_25 (N3708, {N2919, N3450});
or_n #(2, 0, 0) OR_26 (N3709, {N2921, N3451});
or_n #(2, 0, 0) OR_27 (N3710, {N2922, N3452});
or_n #(3, 0, 0) OR_28 (N3711, {N2923, N3453, N503_6});
or_n #(3, 0, 0) OR_29 (N3712, {N2924, N3454, N523_6});
or_n #(3, 0, 0) OR_30 (N3713, {N2925, N3455, N534_6});
or_n #(2, 0, 0) OR_31 (N3715, {N2934, N3459});
or_n #(2, 0, 0) OR_32 (N3716, {N2935, N3460});
or_n #(2, 0, 0) OR_33 (N3717, {N2936, N3461});
or_n #(2, 0, 0) OR_34 (N3718, {N2937, N3462});
or_n #(3, 0, 0) OR_35 (N3719, {N2938, N3463, N389_7});
or_n #(3, 0, 0) OR_36 (N3720, {N2939, N3464, N400_7});
or_n #(3, 0, 0) OR_37 (N3721, {N2940, N3465, N411_7});
or_n #(3, 0, 0) OR_38 (N3722, {N2941, N3466, N374_7});
and_n #(2, 0, 0) AND_260 (N3723, {N369_1, N2942_0});
and_n #(2, 0, 0) AND_261 (N3724, {N361_3, N2942_1});
and_n #(2, 0, 0) AND_262 (N3725, {N351_5, N2942_2});
and_n #(2, 0, 0) AND_263 (N3726, {N341_5, N2942_3});
and_n #(2, 0, 0) AND_264 (N3727, {N324_5, N2948_0});
and_n #(2, 0, 0) AND_265 (N3728, {N316_5, N2948_1});
and_n #(2, 0, 0) AND_266 (N3729, {N308_5, N2948_2});
and_n #(2, 0, 0) AND_267 (N3730, {N302_3, N2948_3});
and_n #(2, 0, 0) AND_268 (N3731, {N293_4, N2948_4});
or_n #(2, 0, 0) OR_39 (N3732, {N2942_4, N2958});
and_n #(2, 0, 0) AND_269 (N3738, {N83_1, N2964_0});
and_n #(2, 0, 0) AND_270 (N3739, {N87, N2964_1});
and_n #(2, 0, 0) AND_271 (N3740, {N34_0, N2964_2});
and_n #(2, 0, 0) AND_272 (N3741, {N34_1, N2964_3});
or_n #(2, 0, 0) OR_40 (N3742, {N2979, N3481});
or_n #(2, 0, 0) OR_41 (N3743, {N2981, N3483});
or_n #(2, 0, 0) OR_42 (N3744, {N2982, N3484});
or_n #(3, 0, 0) OR_43 (N3745, {N2983, N3485, N503_7});
or_n #(3, 0, 0) OR_44 (N3746, {N2985, N3486, N523_7});
or_n #(3, 0, 0) OR_45 (N3747, {N2986, N3487, N534_7});
or_n #(2, 0, 0) OR_46 (N3748, {N2993, N3488});
or_n #(2, 0, 0) OR_47 (N3749, {N2994, N3489});
or_n #(2, 0, 0) OR_48 (N3750, {N2995, N3490});
or_n #(3, 0, 0) OR_49 (N3751, {N2997, N3492, N479_7});
or_n #(3, 0, 0) OR_50 (N3752, {N2998, N3493, N490_7});
notg #(0, 0) NOT_175 (N3753, N3000_0);
notg #(0, 0) NOT_176 (N3754, N3003_0);
notg #(0, 0) NOT_177 (N3755, N3007_0);
notg #(0, 0) NOT_178 (N3756, N3010_0);
or_n #(2, 0, 0) OR_51 (N3757, {N3013, N3502});
and_n #(3, 0, 0) AND_273 (N3758, {N1315_9, N446_2, N3003_1});
or_n #(2, 0, 0) OR_52 (N3759, {N3014, N3503});
and_n #(3, 0, 0) AND_274 (N3760, {N1315_10, N446_3, N3010_1});
and_n #(2, 0, 0) AND_275 (N3761, {N1675_7, N3000_1});
and_n #(2, 0, 0) AND_276 (N3762, {N1675_8, N3007_1});
or_n #(2, 0, 0) OR_53 (N3763, {N3023, N3504});
or_n #(2, 0, 0) OR_54 (N3764, {N3024, N3505});
or_n #(2, 0, 0) OR_55 (N3765, {N3025, N3506});
or_n #(2, 0, 0) OR_56 (N3766, {N3026, N3507});
or_n #(3, 0, 0) OR_57 (N3767, {N3027, N3508, N457_7});
or_n #(3, 0, 0) OR_58 (N3768, {N3028, N3509, N468_7});
or_n #(3, 0, 0) OR_59 (N3769, {N3029, N3510, N422_7});
or_n #(3, 0, 0) OR_60 (N3770, {N3030, N3511, N435_7});
nand_n #(2, 0, 0) NAND_19 (N3771, {N3512, N3513});
nand_n #(2, 0, 0) NAND_20 (N3775, {N3514, N3515});
notg #(0, 0) NOT_179 (N3779, N3035_0);
notg #(0, 0) NOT_180 (N3780, N3038_0);
and_n #(3, 0, 0) AND_277 (N3781, {N117, N3097_1, N1769_3});
and_n #(3, 0, 0) AND_278 (N3782, {N126, N3097_2, N1769_4});
and_n #(3, 0, 0) AND_279 (N3783, {N127, N3097_3, N1769_5});
and_n #(3, 0, 0) AND_280 (N3784, {N128, N3097_4, N1769_6});
and_n #(3, 0, 0) AND_281 (N3785, {N131, N3119_1, N1785_3});
and_n #(3, 0, 0) AND_282 (N3786, {N129, N3119_2, N1785_4});
and_n #(3, 0, 0) AND_283 (N3787, {N119, N3119_3, N1785_5});
and_n #(3, 0, 0) AND_284 (N3788, {N130, N3119_4, N1785_6});
nand_n #(2, 0, 0) NAND_21 (N3789, {N3558, N3559});
nand_n #(2, 0, 0) NAND_22 (N3793, {N3560, N3561});
nand_n #(2, 0, 0) NAND_23 (N3797, {N3562, N3563});
and_n #(3, 0, 0) AND_285 (N3800, {N122, N3147_0, N1800_1});
and_n #(3, 0, 0) AND_286 (N3801, {N113, N3147_1, N1800_2});
and_n #(3, 0, 0) AND_287 (N3802, {N53, N3147_2, N1800_3});
and_n #(3, 0, 0) AND_288 (N3803, {N114, N3147_3, N1800_4});
and_n #(3, 0, 0) AND_289 (N3804, {N115, N3147_4, N1800_5});
and_n #(3, 0, 0) AND_290 (N3805, {N52, N3169_0, N1814_1});
and_n #(3, 0, 0) AND_291 (N3806, {N112, N3169_1, N1814_2});
and_n #(3, 0, 0) AND_292 (N3807, {N116, N3169_2, N1814_3});
and_n #(3, 0, 0) AND_293 (N3808, {N121, N3169_3, N1814_4});
and_n #(3, 0, 0) AND_294 (N3809, {N123_1, N3169_4, N1814_5});
nand_n #(2, 0, 0) NAND_24 (N3810, {N3607, N3608});
nand_n #(2, 0, 0) NAND_25 (N3813, {N3605, N3606});
and_n #(2, 0, 0) AND_295 (N3816, {N3482, N2984});
or_n #(2, 0, 0) OR_61 (N3819, {N2996, N3491});
notg #(0, 0) NOT_181 (N3822, N3200_0);
nand_n #(2, 0, 0) NAND_26 (N3823, {N3200_1, N3203});
nand_n #(2, 0, 0) NAND_27 (N3824, {N3609, N3610});
notg #(0, 0) NOT_182 (N3827, N3456_0);
or_n #(2, 0, 0) OR_62 (N3828, {N3739, N2970});
or_n #(2, 0, 0) OR_63 (N3829, {N3740, N2971});
or_n #(2, 0, 0) OR_64 (N3830, {N3741, N2972});
or_n #(2, 0, 0) OR_65 (N3831, {N3738, N2969});
notg #(0, 0) NOT_183 (N3834, N3664);
notg #(0, 0) NOT_184 (N3835, N3665);
notg #(0, 0) NOT_185 (N3836, N3666);
notg #(0, 0) NOT_186 (N3837, N3667);
notg #(0, 0) NOT_187 (N3838, N3672);
notg #(0, 0) NOT_188 (N3839, N3673);
notg #(0, 0) NOT_189 (N3840, N3674);
notg #(0, 0) NOT_190 (N3841, N3675);
or_n #(2, 0, 0) OR_66 (N3842, {N3681, N2868});
or_n #(2, 0, 0) OR_67 (N3849, {N3682, N2869});
or_n #(2, 0, 0) OR_68 (N3855, {N3683, N2870});
or_n #(2, 0, 0) OR_69 (N3861, {N3684, N2871});
or_n #(2, 0, 0) OR_70 (N3867, {N3685, N2872});
or_n #(2, 0, 0) OR_71 (N3873, {N3686, N2873});
or_n #(2, 0, 0) OR_72 (N3881, {N3687, N2874});
or_n #(2, 0, 0) OR_73 (N3887, {N3688, N2875});
or_n #(2, 0, 0) OR_74 (N3893, {N3689, N2876});
notg #(0, 0) NOT_191 (N3908, N3701);
notg #(0, 0) NOT_192 (N3909, N3702);
notg #(0, 0) NOT_193 (N3911, N3700);
notg #(0, 0) NOT_194 (N3914, N3708);
notg #(0, 0) NOT_195 (N3915, N3709);
notg #(0, 0) NOT_196 (N3916, N3710);
notg #(0, 0) NOT_197 (N3917, N3715);
notg #(0, 0) NOT_198 (N3918, N3716);
notg #(0, 0) NOT_199 (N3919, N3717);
notg #(0, 0) NOT_200 (N3920, N3718);
or_n #(2, 0, 0) OR_75 (N3921, {N3724, N2955});
or_n #(2, 0, 0) OR_76 (N3927, {N3725, N2956});
or_n #(2, 0, 0) OR_77 (N3933, {N3726, N2957});
or_n #(2, 0, 0) OR_78 (N3942, {N3727, N2959});
or_n #(2, 0, 0) OR_79 (N3948, {N3728, N2960});
or_n #(2, 0, 0) OR_80 (N3956, {N3729, N2961});
or_n #(2, 0, 0) OR_81 (N3962, {N3730, N2962});
or_n #(2, 0, 0) OR_82 (N3968, {N3731, N2963});
notg #(0, 0) NOT_201 (N3975, N3742);
notg #(0, 0) NOT_202 (N3976, N3743);
notg #(0, 0) NOT_203 (N3977, N3744);
notg #(0, 0) NOT_204 (N3978, N3749);
notg #(0, 0) NOT_205 (N3979, N3750);
and_n #(3, 0, 0) AND_296 (N3980, {N446_4, N1292_8, N3754});
and_n #(3, 0, 0) AND_297 (N3981, {N446_5, N1292_9, N3756});
and_n #(2, 0, 0) AND_298 (N3982, {N1271_6, N3753});
and_n #(2, 0, 0) AND_299 (N3983, {N1271_7, N3755});
notg #(0, 0) NOT_206 (N3984, N3757);
notg #(0, 0) NOT_207 (N3987, N3759);
notg #(0, 0) NOT_208 (N3988, N3763);
notg #(0, 0) NOT_209 (N3989, N3764);
notg #(0, 0) NOT_210 (N3990, N3765);
notg #(0, 0) NOT_211 (N3991, N3766);
and_n #(3, 0, 0) AND_300 (N3998, {N3456_1, N3119_5, N3130_0});
or_n #(2, 0, 0) OR_83 (N4008, {N3723, N2954});
or_n #(2, 0, 0) OR_84 (N4011, {N3680, N2867});
notg #(0, 0) NOT_212 (N4021, N3748);
nand_n #(2, 0, 0) NAND_28 (N4024, {N1968_1, N3822});
notg #(0, 0) NOT_213 (N4027, N3705_0);
and_n #(2, 0, 0) AND_301 (N4031, {N3828, N1583_0});
and_n #(3, 0, 0) AND_302 (N4032, {N24, N2882_4, N3691_0});
and_n #(3, 0, 0) AND_303 (N4033, {N25, N1482_5, N3691_1});
and_n #(3, 0, 0) AND_304 (N4034, {N26, N2882_5, N3691_2});
and_n #(3, 0, 0) AND_305 (N4035, {N81, N1482_6, N3691_3});
and_n #(2, 0, 0) AND_306 (N4036, {N3829, N1583_1});
and_n #(3, 0, 0) AND_307 (N4037, {N79, N2882_6, N3691_4});
and_n #(3, 0, 0) AND_308 (N4038, {N23, N1482_7, N3691_5});
and_n #(3, 0, 0) AND_309 (N4039, {N82, N2882_7, N3691_6});
and_n #(3, 0, 0) AND_310 (N4040, {N80, N1482_8, N3691_7});
and_n #(2, 0, 0) AND_311 (N4041, {N3830, N1583_2});
and_n #(2, 0, 0) AND_312 (N4042, {N3831, N1583_3});
and_n #(2, 0, 0) AND_313 (N4067, {N3732_0, N514_6});
and_n #(2, 0, 0) AND_314 (N4080, {N514_7, N3732_1});
and_n #(2, 0, 0) AND_315 (N4088, {N3834, N3668});
and_n #(2, 0, 0) AND_316 (N4091, {N3835, N3669});
and_n #(2, 0, 0) AND_317 (N4094, {N3836, N3670});
and_n #(2, 0, 0) AND_318 (N4097, {N3837, N3671});
and_n #(2, 0, 0) AND_319 (N4100, {N3838, N3676});
and_n #(2, 0, 0) AND_320 (N4103, {N3839, N3677});
and_n #(2, 0, 0) AND_321 (N4106, {N3840, N3678});
and_n #(2, 0, 0) AND_322 (N4109, {N3841, N3679});
and_n #(2, 0, 0) AND_323 (N4144, {N3908, N3703});
and_n #(2, 0, 0) AND_324 (N4147, {N3909, N3704});
bufg #(0, 0) BUF_181 (N4150, N3705_1);
and_n #(2, 0, 0) AND_325 (N4153, {N3914, N3711});
and_n #(2, 0, 0) AND_326 (N4156, {N3915, N3712});
and_n #(2, 0, 0) AND_327 (N4159, {N3916, N3713});
or_n #(2, 0, 0) OR_85 (N4183, {N3758, N3980});
or_n #(2, 0, 0) OR_86 (N4184, {N3760, N3981});
or_n #(3, 0, 0) OR_87 (N4185, {N3761, N3982, N446_6});
or_n #(3, 0, 0) OR_88 (N4186, {N3762, N3983, N446_7});
notg #(0, 0) NOT_214 (N4188, N3771_0);
notg #(0, 0) NOT_215 (N4191, N3775_0);
and_n #(3, 0, 0) AND_328 (N4196, {N3775_1, N3771_1, N3035_1});
and_n #(3, 0, 0) AND_329 (N4197, {N3987, N3119_6, N3130_1});
and_n #(2, 0, 0) AND_330 (N4198, {N3920, N3722});
notg #(0, 0) NOT_216 (N4199, N3816_0);
notg #(0, 0) NOT_217 (N4200, N3789_0);
notg #(0, 0) NOT_218 (N4203, N3793_0);
bufg #(0, 0) BUF_182 (N4206, N3797_0);
bufg #(0, 0) BUF_183 (N4209, N3797_1);
bufg #(0, 0) BUF_184 (N4212, N3732_2);
bufg #(0, 0) BUF_185 (N4215, N3732_3);
bufg #(0, 0) BUF_186 (N4219, N3732_4);
notg #(0, 0) NOT_219 (N4223, N3810_0);
notg #(0, 0) NOT_220 (N4224, N3813_0);
and_n #(2, 0, 0) AND_331 (N4225, {N3918, N3720});
and_n #(2, 0, 0) AND_332 (N4228, {N3919, N3721});
and_n #(2, 0, 0) AND_333 (N4231, {N3991, N3770});
and_n #(2, 0, 0) AND_334 (N4234, {N3917, N3719});
and_n #(2, 0, 0) AND_335 (N4237, {N3989, N3768});
and_n #(2, 0, 0) AND_336 (N4240, {N3990, N3769});
and_n #(2, 0, 0) AND_337 (N4243, {N3988, N3767});
and_n #(2, 0, 0) AND_338 (N4246, {N3976, N3746});
and_n #(2, 0, 0) AND_339 (N4249, {N3977, N3747});
and_n #(2, 0, 0) AND_340 (N4252, {N3975, N3745});
and_n #(2, 0, 0) AND_341 (N4255, {N3978, N3751});
and_n #(2, 0, 0) AND_342 (N4258, {N3979, N3752});
notg #(0, 0) NOT_221 (N4263, N3819_0);
nand_n #(2, 0, 0) NAND_29 (N4264, {N4024, N3823});
notg #(0, 0) NOT_222 (N4267, N3824_0);
and_n #(2, 0, 0) AND_343 (N4268, {N446_8, N3893_0});
notg #(0, 0) NOT_223 (N4269, N3911_0);
notg #(0, 0) NOT_224 (N4270, N3984_0);
and_n #(2, 0, 0) AND_344 (N4271, {N3893_1, N446_9});
notg #(0, 0) NOT_225 (N4272, N4031);
or_n #(4, 0, 0) OR_89 (N4273, {N4032, N4033, N3614, N3615});
or_n #(4, 0, 0) OR_90 (N4274, {N4034, N4035, N3625, N3626});
notg #(0, 0) NOT_226 (N4275, N4036);
or_n #(4, 0, 0) OR_91 (N4276, {N4037, N4038, N3636, N3637});
or_n #(4, 0, 0) OR_92 (N4277, {N4039, N4040, N3639, N3640});
notg #(0, 0) NOT_227 (N4278, N4041);
notg #(0, 0) NOT_228 (N4279, N4042);
and_n #(2, 0, 0) AND_345 (N4280, {N3887_0, N457_8});
and_n #(2, 0, 0) AND_346 (N4284, {N3881_0, N468_8});
and_n #(2, 0, 0) AND_347 (N4290, {N422_8, N3873_0});
and_n #(2, 0, 0) AND_348 (N4297, {N3867_0, N435_8});
and_n #(2, 0, 0) AND_349 (N4298, {N3861_0, N389_8});
and_n #(2, 0, 0) AND_350 (N4301, {N3855_0, N400_8});
and_n #(2, 0, 0) AND_351 (N4305, {N3849_0, N411_8});
and_n #(2, 0, 0) AND_352 (N4310, {N3842_0, N374_8});
and_n #(2, 0, 0) AND_353 (N4316, {N457_9, N3887_1});
and_n #(2, 0, 0) AND_354 (N4320, {N468_9, N3881_1});
and_n #(2, 0, 0) AND_355 (N4325, {N422_9, N3873_1});
and_n #(2, 0, 0) AND_356 (N4331, {N435_9, N3867_1});
and_n #(2, 0, 0) AND_357 (N4332, {N389_9, N3861_1});
and_n #(2, 0, 0) AND_358 (N4336, {N400_9, N3855_1});
and_n #(2, 0, 0) AND_359 (N4342, {N411_9, N3849_1});
and_n #(2, 0, 0) AND_360 (N4349, {N374_9, N3842_1});
notg #(0, 0) NOT_229 (N4357, N3968_0);
notg #(0, 0) NOT_230 (N4364, N3962_0);
bufg #(0, 0) BUF_187 (N4375, N3962_1);
and_n #(2, 0, 0) AND_361 (N4379, {N3956_0, N479_8});
and_n #(2, 0, 0) AND_362 (N4385, {N490_8, N3948_0});
and_n #(2, 0, 0) AND_363 (N4392, {N3942_0, N503_8});
and_n #(2, 0, 0) AND_364 (N4396, {N3933_0, N523_8});
and_n #(2, 0, 0) AND_365 (N4400, {N3927_0, N534_8});
notg #(0, 0) NOT_231 (N4405, N3921_0);
bufg #(0, 0) BUF_188 (N4412, N3921_1);
notg #(0, 0) NOT_232 (N4418, N3968_1);
notg #(0, 0) NOT_233 (N4425, N3962_2);
bufg #(0, 0) BUF_189 (N4436, N3962_3);
and_n #(2, 0, 0) AND_366 (N4440, {N479_9, N3956_1});
and_n #(2, 0, 0) AND_367 (N4445, {N490_9, N3948_1});
and_n #(2, 0, 0) AND_368 (N4451, {N503_9, N3942_1});
and_n #(2, 0, 0) AND_369 (N4456, {N523_9, N3933_1});
and_n #(2, 0, 0) AND_370 (N4462, {N534_9, N3927_1});
bufg #(0, 0) BUF_190 (N4469, N3921_2);
notg #(0, 0) NOT_234 (N4477, N3921_3);
bufg #(0, 0) BUF_191 (N4512, N3968_2);
notg #(0, 0) NOT_235 (N4515, N4183);
notg #(0, 0) NOT_236 (N4516, N4184);
notg #(0, 0) NOT_237 (N4521, N4008_0);
notg #(0, 0) NOT_238 (N4523, N4011_0);
notg #(0, 0) NOT_239 (N4524, N4198);
notg #(0, 0) NOT_240 (N4532, N3984_1);
and_n #(3, 0, 0) AND_371 (N4547, {N3911_1, N3169_5, N3180_0});
bufg #(0, 0) BUF_192 (N4548, N3893_2);
bufg #(0, 0) BUF_193 (N4551, N3887_2);
bufg #(0, 0) BUF_194 (N4554, N3881_2);
bufg #(0, 0) BUF_195 (N4557, N3873_2);
bufg #(0, 0) BUF_196 (N4560, N3867_2);
bufg #(0, 0) BUF_197 (N4563, N3861_2);
bufg #(0, 0) BUF_198 (N4566, N3855_2);
bufg #(0, 0) BUF_199 (N4569, N3849_2);
bufg #(0, 0) BUF_200 (N4572, N3842_2);
nor_n #(2, 0, 0) NOR_1 (N4575, {N422_10, N3873_3});
bufg #(0, 0) BUF_201 (N4578, N3893_3);
bufg #(0, 0) BUF_202 (N4581, N3887_3);
bufg #(0, 0) BUF_203 (N4584, N3881_3);
bufg #(0, 0) BUF_204 (N4587, N3867_3);
bufg #(0, 0) BUF_205 (N4590, N3861_3);
bufg #(0, 0) BUF_206 (N4593, N3855_3);
bufg #(0, 0) BUF_207 (N4596, N3849_3);
bufg #(0, 0) BUF_208 (N4599, N3873_4);
bufg #(0, 0) BUF_209 (N4602, N3842_3);
nor_n #(2, 0, 0) NOR_2 (N4605, {N422_11, N3873_5});
nor_n #(2, 0, 0) NOR_3 (N4608, {N374_10, N3842_4});
bufg #(0, 0) BUF_210 (N4611, N3956_2);
bufg #(0, 0) BUF_211 (N4614, N3948_2);
bufg #(0, 0) BUF_212 (N4617, N3942_2);
bufg #(0, 0) BUF_213 (N4621, N3933_2);
bufg #(0, 0) BUF_214 (N4624, N3927_2);
nor_n #(2, 0, 0) NOR_4 (N4627, {N490_10, N3948_3});
bufg #(0, 0) BUF_215 (N4630, N3956_3);
bufg #(0, 0) BUF_216 (N4633, N3942_3);
bufg #(0, 0) BUF_217 (N4637, N3933_3);
bufg #(0, 0) BUF_218 (N4640, N3927_3);
bufg #(0, 0) BUF_219 (N4643, N3948_4);
nor_n #(2, 0, 0) NOR_5 (N4646, {N490_11, N3948_5});
bufg #(0, 0) BUF_220 (N4649, N3927_4);
bufg #(0, 0) BUF_221 (N4652, N3933_4);
bufg #(0, 0) BUF_222 (N4655, N3921_4);
bufg #(0, 0) BUF_223 (N4658, N3942_4);
bufg #(0, 0) BUF_224 (N4662, N3956_4);
bufg #(0, 0) BUF_225 (N4665, N3948_6);
bufg #(0, 0) BUF_226 (N4668, N3968_3);
bufg #(0, 0) BUF_227 (N4671, N3962_4);
bufg #(0, 0) BUF_228 (N4674, N3873_6);
bufg #(0, 0) BUF_229 (N4677, N3867_4);
bufg #(0, 0) BUF_230 (N4680, N3887_4);
bufg #(0, 0) BUF_231 (N4683, N3881_4);
bufg #(0, 0) BUF_232 (N4686, N3893_4);
bufg #(0, 0) BUF_233 (N4689, N3849_4);
bufg #(0, 0) BUF_234 (N4692, N3842_5);
bufg #(0, 0) BUF_235 (N4695, N3861_4);
bufg #(0, 0) BUF_236 (N4698, N3855_4);
nand_n #(2, 0, 0) NAND_30 (N4701, {N3813_1, N4223});
nand_n #(2, 0, 0) NAND_31 (N4702, {N3810_1, N4224});
notg #(0, 0) NOT_241 (N4720, N4021_0);
nand_n #(2, 0, 0) NAND_32 (N4721, {N4021_1, N4263});
notg #(0, 0) NOT_242 (N4724, N4147_0);
notg #(0, 0) NOT_243 (N4725, N4144_0);
notg #(0, 0) NOT_244 (N4726, N4159_0);
notg #(0, 0) NOT_245 (N4727, N4156_0);
notg #(0, 0) NOT_246 (N4728, N4153_0);
notg #(0, 0) NOT_247 (N4729, N4097_0);
notg #(0, 0) NOT_248 (N4730, N4094_0);
notg #(0, 0) NOT_249 (N4731, N4091_0);
notg #(0, 0) NOT_250 (N4732, N4088_0);
notg #(0, 0) NOT_251 (N4733, N4109_0);
notg #(0, 0) NOT_252 (N4734, N4106_0);
notg #(0, 0) NOT_253 (N4735, N4103_0);
notg #(0, 0) NOT_254 (N4736, N4100_0);
and_n #(2, 0, 0) AND_372 (N4737, {N4273, N2877_0});
and_n #(2, 0, 0) AND_373 (N4738, {N4274, N2877_1});
and_n #(2, 0, 0) AND_374 (N4739, {N4276, N2877_2});
and_n #(2, 0, 0) AND_375 (N4740, {N4277, N2877_3});
and_n #(3, 0, 0) AND_376 (N4741, {N4150_0, N1758_1, N1755_0});
notg #(0, 0) NOT_255 (N4855, N4212_0);
nand_n #(2, 0, 0) NAND_33 (N4856, {N4212_1, N2712});
nand_n #(2, 0, 0) NAND_34 (N4908, {N4215_0, N2718});
notg #(0, 0) NOT_256 (N4909, N4215_1);
and_n #(2, 0, 0) AND_377 (N4939, {N4515, N4185});
and_n #(2, 0, 0) AND_378 (N4942, {N4516, N4186});
notg #(0, 0) NOT_257 (N4947, N4219_0);
and_n #(3, 0, 0) AND_379 (N4953, {N4188_0, N3775_2, N3779});
and_n #(3, 0, 0) AND_380 (N4954, {N3771_2, N4191_0, N3780});
and_n #(3, 0, 0) AND_381 (N4955, {N4191_1, N4188_1, N3038_1});
and_n #(3, 0, 0) AND_382 (N4956, {N4109_1, N3097_5, N3108_0});
and_n #(3, 0, 0) AND_383 (N4957, {N4106_1, N3097_6, N3108_1});
and_n #(3, 0, 0) AND_384 (N4958, {N4103_1, N3097_7, N3108_2});
and_n #(3, 0, 0) AND_385 (N4959, {N4100_1, N3097_8, N3108_3});
and_n #(3, 0, 0) AND_386 (N4960, {N4159_1, N3119_7, N3130_2});
and_n #(3, 0, 0) AND_387 (N4961, {N4156_1, N3119_8, N3130_3});
notg #(0, 0) NOT_258 (N4965, N4225_0);
notg #(0, 0) NOT_259 (N4966, N4228_0);
notg #(0, 0) NOT_260 (N4967, N4231_0);
notg #(0, 0) NOT_261 (N4968, N4234_0);
notg #(0, 0) NOT_262 (N4972, N4246_0);
notg #(0, 0) NOT_263 (N4973, N4249_0);
notg #(0, 0) NOT_264 (N4974, N4252_0);
nand_n #(2, 0, 0) NAND_35 (N4975, {N4252_1, N4199});
notg #(0, 0) NOT_265 (N4976, N4206_0);
notg #(0, 0) NOT_266 (N4977, N4209_0);
and_n #(3, 0, 0) AND_388 (N4978, {N3793_1, N3789_1, N4206_1});
and_n #(3, 0, 0) AND_389 (N4979, {N4203_0, N4200_0, N4209_1});
and_n #(3, 0, 0) AND_390 (N4980, {N4097_1, N3147_5, N3158_0});
and_n #(3, 0, 0) AND_391 (N4981, {N4094_1, N3147_6, N3158_1});
and_n #(3, 0, 0) AND_392 (N4982, {N4091_1, N3147_7, N3158_2});
and_n #(3, 0, 0) AND_393 (N4983, {N4088_1, N3147_8, N3158_3});
and_n #(3, 0, 0) AND_394 (N4984, {N4153_1, N3169_6, N3180_1});
and_n #(3, 0, 0) AND_395 (N4985, {N4147_1, N3169_7, N3180_2});
and_n #(3, 0, 0) AND_396 (N4986, {N4144_1, N3169_8, N3180_3});
and_n #(3, 0, 0) AND_397 (N4987, {N4150_1, N3169_9, N3180_4});
nand_n #(2, 0, 0) NAND_36 (N5049, {N4701, N4702});
notg #(0, 0) NOT_267 (N5052, N4237_0);
notg #(0, 0) NOT_268 (N5053, N4240_0);
notg #(0, 0) NOT_269 (N5054, N4243_0);
notg #(0, 0) NOT_270 (N5055, N4255_0);
notg #(0, 0) NOT_271 (N5056, N4258_0);
nand_n #(2, 0, 0) NAND_37 (N5057, {N3819_1, N4720});
notg #(0, 0) NOT_272 (N5058, N4264_0);
nand_n #(2, 0, 0) NAND_38 (N5059, {N4264_1, N4267});
and_n #(4, 0, 0) AND_398 (N5060, {N4724, N4725, N4269, N4027});
and_n #(4, 0, 0) AND_399 (N5061, {N4726, N4727, N3827, N4728});
and_n #(4, 0, 0) AND_400 (N5062, {N4729, N4730, N4731, N4732});
and_n #(4, 0, 0) AND_401 (N5063, {N4733, N4734, N4735, N4736});
and_n #(2, 0, 0) AND_402 (N5065, {N4357_0, N4375_0});
and_n #(3, 0, 0) AND_403 (N5066, {N4364_0, N4357_1, N4379_0});
and_n #(2, 0, 0) AND_404 (N5067, {N4418_0, N4436_0});
and_n #(3, 0, 0) AND_405 (N5068, {N4425_0, N4418_1, N4440_0});
notg #(0, 0) NOT_273 (N5069, N4548_0);
nand_n #(2, 0, 0) NAND_39 (N5070, {N4548_1, N2628});
notg #(0, 0) NOT_274 (N5071, N4551_0);
nand_n #(2, 0, 0) NAND_40 (N5072, {N4551_1, N2629});
notg #(0, 0) NOT_275 (N5073, N4554_0);
nand_n #(2, 0, 0) NAND_41 (N5074, {N4554_1, N2630});
notg #(0, 0) NOT_276 (N5075, N4557_0);
nand_n #(2, 0, 0) NAND_42 (N5076, {N4557_1, N2631});
notg #(0, 0) NOT_277 (N5077, N4560_0);
nand_n #(2, 0, 0) NAND_43 (N5078, {N4560_1, N2632});
notg #(0, 0) NOT_278 (N5079, N4563_0);
nand_n #(2, 0, 0) NAND_44 (N5080, {N4563_1, N2633});
notg #(0, 0) NOT_279 (N5081, N4566_0);
nand_n #(2, 0, 0) NAND_45 (N5082, {N4566_1, N2634});
notg #(0, 0) NOT_280 (N5083, N4569_0);
nand_n #(2, 0, 0) NAND_46 (N5084, {N4569_1, N2635});
notg #(0, 0) NOT_281 (N5085, N4572_0);
nand_n #(2, 0, 0) NAND_47 (N5086, {N4572_1, N2636});
notg #(0, 0) NOT_282 (N5087, N4575_0);
nand_n #(2, 0, 0) NAND_48 (N5088, {N4578_0, N2638});
notg #(0, 0) NOT_283 (N5089, N4578_1);
nand_n #(2, 0, 0) NAND_49 (N5090, {N4581_0, N2639});
notg #(0, 0) NOT_284 (N5091, N4581_1);
nand_n #(2, 0, 0) NAND_50 (N5092, {N4584_0, N2640});
notg #(0, 0) NOT_285 (N5093, N4584_1);
nand_n #(2, 0, 0) NAND_51 (N5094, {N4587_0, N2641});
notg #(0, 0) NOT_286 (N5095, N4587_1);
nand_n #(2, 0, 0) NAND_52 (N5096, {N4590_0, N2642});
notg #(0, 0) NOT_287 (N5097, N4590_1);
nand_n #(2, 0, 0) NAND_53 (N5098, {N4593_0, N2643});
notg #(0, 0) NOT_288 (N5099, N4593_1);
nand_n #(2, 0, 0) NAND_54 (N5100, {N4596_0, N2644});
notg #(0, 0) NOT_289 (N5101, N4596_1);
nand_n #(2, 0, 0) NAND_55 (N5102, {N4599_0, N2645});
notg #(0, 0) NOT_290 (N5103, N4599_1);
nand_n #(2, 0, 0) NAND_56 (N5104, {N4602_0, N2646});
notg #(0, 0) NOT_291 (N5105, N4602_1);
notg #(0, 0) NOT_292 (N5106, N4611_0);
nand_n #(2, 0, 0) NAND_57 (N5107, {N4611_1, N2709});
notg #(0, 0) NOT_293 (N5108, N4614_0);
nand_n #(2, 0, 0) NAND_58 (N5109, {N4614_1, N2710});
notg #(0, 0) NOT_294 (N5110, N4617_0);
nand_n #(2, 0, 0) NAND_59 (N5111, {N4617_1, N2711});
nand_n #(2, 0, 0) NAND_60 (N5112, {N1890_1, N4855});
notg #(0, 0) NOT_295 (N5113, N4621_0);
nand_n #(2, 0, 0) NAND_61 (N5114, {N4621_1, N2713});
notg #(0, 0) NOT_296 (N5115, N4624_0);
nand_n #(2, 0, 0) NAND_62 (N5116, {N4624_1, N2714});
and_n #(2, 0, 0) AND_406 (N5117, {N4364_1, N4379_1});
and_n #(2, 0, 0) AND_407 (N5118, {N4364_2, N4379_2});
and_n #(2, 0, 0) AND_408 (N5119, {N54_1, N4405_0});
notg #(0, 0) NOT_297 (N5120, N4627_0);
nand_n #(2, 0, 0) NAND_63 (N5121, {N4630_0, N2716});
notg #(0, 0) NOT_298 (N5122, N4630_1);
nand_n #(2, 0, 0) NAND_64 (N5123, {N4633_0, N2717});
notg #(0, 0) NOT_299 (N5124, N4633_1);
nand_n #(2, 0, 0) NAND_65 (N5125, {N1908_1, N4909});
nand_n #(2, 0, 0) NAND_66 (N5126, {N4637_0, N2719});
notg #(0, 0) NOT_300 (N5127, N4637_1);
nand_n #(2, 0, 0) NAND_67 (N5128, {N4640_0, N2720});
notg #(0, 0) NOT_301 (N5129, N4640_1);
nand_n #(2, 0, 0) NAND_68 (N5130, {N4643_0, N2721});
notg #(0, 0) NOT_302 (N5131, N4643_1);
and_n #(2, 0, 0) AND_409 (N5132, {N4425_1, N4440_1});
and_n #(2, 0, 0) AND_410 (N5133, {N4425_2, N4440_2});
notg #(0, 0) NOT_303 (N5135, N4649_0);
notg #(0, 0) NOT_304 (N5136, N4652_0);
nand_n #(2, 0, 0) NAND_69 (N5137, {N4655_0, N4521});
notg #(0, 0) NOT_305 (N5138, N4655_1);
notg #(0, 0) NOT_306 (N5139, N4658_0);
nand_n #(2, 0, 0) NAND_70 (N5140, {N4658_1, N4947});
notg #(0, 0) NOT_307 (N5141, N4674_0);
notg #(0, 0) NOT_308 (N5142, N4677_0);
notg #(0, 0) NOT_309 (N5143, N4680_0);
notg #(0, 0) NOT_310 (N5144, N4683_0);
nand_n #(2, 0, 0) NAND_71 (N5145, {N4686_0, N4523});
notg #(0, 0) NOT_311 (N5146, N4686_1);
nor_n #(2, 0, 0) NOR_6 (N5147, {N4953, N4196});
nor_n #(2, 0, 0) NOR_7 (N5148, {N4954, N4955});
notg #(0, 0) NOT_312 (N5150, N4524_0);
nand_n #(2, 0, 0) NAND_72 (N5153, {N4228_1, N4965});
nand_n #(2, 0, 0) NAND_73 (N5154, {N4225_1, N4966});
nand_n #(2, 0, 0) NAND_74 (N5155, {N4234_1, N4967});
nand_n #(2, 0, 0) NAND_75 (N5156, {N4231_1, N4968});
notg #(0, 0) NOT_313 (N5157, N4532_0);
nand_n #(2, 0, 0) NAND_76 (N5160, {N4249_1, N4972});
nand_n #(2, 0, 0) NAND_77 (N5161, {N4246_1, N4973});
nand_n #(2, 0, 0) NAND_78 (N5162, {N3816_1, N4974});
and_n #(3, 0, 0) AND_411 (N5163, {N4200_1, N3793_2, N4976});
and_n #(3, 0, 0) AND_412 (N5164, {N3789_2, N4203_1, N4977});
and_n #(3, 0, 0) AND_413 (N5165, {N4942, N3147_9, N3158_4});
notg #(0, 0) NOT_314 (N5166, N4512_0);
bufg #(0, 0) BUF_237 (N5169, N4290_0);
notg #(0, 0) NOT_315 (N5172, N4605_0);
bufg #(0, 0) BUF_238 (N5173, N4325_0);
notg #(0, 0) NOT_316 (N5176, N4608_0);
bufg #(0, 0) BUF_239 (N5177, N4349_0);
bufg #(0, 0) BUF_240 (N5180, N4405_1);
bufg #(0, 0) BUF_241 (N5183, N4357_2);
bufg #(0, 0) BUF_242 (N5186, N4357_3);
bufg #(0, 0) BUF_243 (N5189, N4364_3);
bufg #(0, 0) BUF_244 (N5192, N4364_4);
bufg #(0, 0) BUF_245 (N5195, N4385_0);
notg #(0, 0) NOT_317 (N5198, N4646_0);
bufg #(0, 0) BUF_246 (N5199, N4418_2);
bufg #(0, 0) BUF_247 (N5202, N4425_3);
bufg #(0, 0) BUF_248 (N5205, N4445_0);
bufg #(0, 0) BUF_249 (N5208, N4418_3);
bufg #(0, 0) BUF_250 (N5211, N4425_4);
bufg #(0, 0) BUF_251 (N5214, N4477_0);
bufg #(0, 0) BUF_252 (N5217, N4469_0);
bufg #(0, 0) BUF_253 (N5220, N4477_1);
notg #(0, 0) NOT_318 (N5223, N4662_0);
notg #(0, 0) NOT_319 (N5224, N4665_0);
notg #(0, 0) NOT_320 (N5225, N4668_0);
notg #(0, 0) NOT_321 (N5226, N4671_0);
notg #(0, 0) NOT_322 (N5227, N4689_0);
notg #(0, 0) NOT_323 (N5228, N4692_0);
notg #(0, 0) NOT_324 (N5229, N4695_0);
notg #(0, 0) NOT_325 (N5230, N4698_0);
nand_n #(2, 0, 0) NAND_79 (N5232, {N4240_1, N5052});
nand_n #(2, 0, 0) NAND_80 (N5233, {N4237_1, N5053});
nand_n #(2, 0, 0) NAND_81 (N5234, {N4258_1, N5055});
nand_n #(2, 0, 0) NAND_82 (N5235, {N4255_1, N5056});
nand_n #(2, 0, 0) NAND_83 (N5236, {N4721, N5057});
nand_n #(2, 0, 0) NAND_84 (N5239, {N3824_1, N5058});
and_n #(3, 0, 0) AND_414 (N5240, {N5060, N5061, N4270});
notg #(0, 0) NOT_326 (N5241, N4939_0);
nand_n #(2, 0, 0) NAND_85 (N5242, {N1824_1, N5069});
nand_n #(2, 0, 0) NAND_86 (N5243, {N1827_1, N5071});
nand_n #(2, 0, 0) NAND_87 (N5244, {N1830_1, N5073});
nand_n #(2, 0, 0) NAND_88 (N5245, {N1833_1, N5075});
nand_n #(2, 0, 0) NAND_89 (N5246, {N1836_1, N5077});
nand_n #(2, 0, 0) NAND_90 (N5247, {N1839_1, N5079});
nand_n #(2, 0, 0) NAND_91 (N5248, {N1842_1, N5081});
nand_n #(2, 0, 0) NAND_92 (N5249, {N1845_1, N5083});
nand_n #(2, 0, 0) NAND_93 (N5250, {N1848_1, N5085});
nand_n #(2, 0, 0) NAND_94 (N5252, {N1854_1, N5089});
nand_n #(2, 0, 0) NAND_95 (N5253, {N1857_1, N5091});
nand_n #(2, 0, 0) NAND_96 (N5254, {N1860_1, N5093});
nand_n #(2, 0, 0) NAND_97 (N5255, {N1863_1, N5095});
nand_n #(2, 0, 0) NAND_98 (N5256, {N1866_1, N5097});
nand_n #(2, 0, 0) NAND_99 (N5257, {N1869_1, N5099});
nand_n #(2, 0, 0) NAND_100 (N5258, {N1872_1, N5101});
nand_n #(2, 0, 0) NAND_101 (N5259, {N1875_1, N5103});
nand_n #(2, 0, 0) NAND_102 (N5260, {N1878_1, N5105});
nand_n #(2, 0, 0) NAND_103 (N5261, {N1881_1, N5106});
nand_n #(2, 0, 0) NAND_104 (N5262, {N1884_1, N5108});
nand_n #(2, 0, 0) NAND_105 (N5263, {N1887_1, N5110});
nand_n #(2, 0, 0) NAND_106 (N5264, {N5112, N4856});
nand_n #(2, 0, 0) NAND_107 (N5274, {N1893_1, N5113});
nand_n #(2, 0, 0) NAND_108 (N5275, {N1896_1, N5115});
nand_n #(2, 0, 0) NAND_109 (N5282, {N1902_1, N5122});
nand_n #(2, 0, 0) NAND_110 (N5283, {N1905_1, N5124});
nand_n #(2, 0, 0) NAND_111 (N5284, {N4908, N5125});
nand_n #(2, 0, 0) NAND_112 (N5298, {N1911_1, N5127});
nand_n #(2, 0, 0) NAND_113 (N5299, {N1914_1, N5129});
nand_n #(2, 0, 0) NAND_114 (N5300, {N1917_1, N5131});
nand_n #(2, 0, 0) NAND_115 (N5303, {N4652_1, N5135});
nand_n #(2, 0, 0) NAND_116 (N5304, {N4649_1, N5136});
nand_n #(2, 0, 0) NAND_117 (N5305, {N4008_1, N5138});
nand_n #(2, 0, 0) NAND_118 (N5306, {N4219_1, N5139});
nand_n #(2, 0, 0) NAND_119 (N5307, {N4677_1, N5141});
nand_n #(2, 0, 0) NAND_120 (N5308, {N4674_1, N5142});
nand_n #(2, 0, 0) NAND_121 (N5309, {N4683_1, N5143});
nand_n #(2, 0, 0) NAND_122 (N5310, {N4680_1, N5144});
nand_n #(2, 0, 0) NAND_123 (N5311, {N4011_1, N5146});
notg #(0, 0) NOT_327 (N5312, N5049_0);
nand_n #(2, 0, 0) NAND_124 (N5315, {N5153, N5154});
nand_n #(2, 0, 0) NAND_125 (N5319, {N5155, N5156});
nand_n #(2, 0, 0) NAND_126 (N5324, {N5160, N5161});
nand_n #(2, 0, 0) NAND_127 (N5328, {N5162, N4975});
nor_n #(2, 0, 0) NOR_8 (N5331, {N5163, N4978});
nor_n #(2, 0, 0) NOR_9 (N5332, {N5164, N4979});
or_n #(2, 0, 0) OR_93 (N5346, {N4412_0, N5119});
nand_n #(2, 0, 0) NAND_128 (N5363, {N4665_1, N5223});
nand_n #(2, 0, 0) NAND_129 (N5364, {N4662_1, N5224});
nand_n #(2, 0, 0) NAND_130 (N5365, {N4671_1, N5225});
nand_n #(2, 0, 0) NAND_131 (N5366, {N4668_1, N5226});
nand_n #(2, 0, 0) NAND_132 (N5367, {N4692_1, N5227});
nand_n #(2, 0, 0) NAND_133 (N5368, {N4689_1, N5228});
nand_n #(2, 0, 0) NAND_134 (N5369, {N4698_1, N5229});
nand_n #(2, 0, 0) NAND_135 (N5370, {N4695_1, N5230});
nand_n #(2, 0, 0) NAND_136 (N5371, {N5148, N5147});
bufg #(0, 0) BUF_254 (N5374, N4939_1);
nand_n #(2, 0, 0) NAND_137 (N5377, {N5232, N5233});
nand_n #(2, 0, 0) NAND_138 (N5382, {N5234, N5235});
nand_n #(2, 0, 0) NAND_139 (N5385, {N5239, N5059});
and_n #(3, 0, 0) AND_415 (N5388, {N5062, N5063, N5241});
nand_n #(2, 0, 0) NAND_140 (N5389, {N5242, N5070});
nand_n #(2, 0, 0) NAND_141 (N5396, {N5243, N5072});
nand_n #(2, 0, 0) NAND_142 (N5407, {N5244, N5074});
nand_n #(2, 0, 0) NAND_143 (N5418, {N5245, N5076});
nand_n #(2, 0, 0) NAND_144 (N5424, {N5246, N5078});
nand_n #(2, 0, 0) NAND_145 (N5431, {N5247, N5080});
nand_n #(2, 0, 0) NAND_146 (N5441, {N5248, N5082});
nand_n #(2, 0, 0) NAND_147 (N5452, {N5249, N5084});
nand_n #(2, 0, 0) NAND_148 (N5462, {N5250, N5086});
notg #(0, 0) NOT_328 (N5469, N5169_0);
nand_n #(2, 0, 0) NAND_149 (N5470, {N5088, N5252});
nand_n #(2, 0, 0) NAND_150 (N5477, {N5090, N5253});
nand_n #(2, 0, 0) NAND_151 (N5488, {N5092, N5254});
nand_n #(2, 0, 0) NAND_152 (N5498, {N5094, N5255});
nand_n #(2, 0, 0) NAND_153 (N5506, {N5096, N5256});
nand_n #(2, 0, 0) NAND_154 (N5520, {N5098, N5257});
nand_n #(2, 0, 0) NAND_155 (N5536, {N5100, N5258});
nand_n #(2, 0, 0) NAND_156 (N5549, {N5102, N5259});
nand_n #(2, 0, 0) NAND_157 (N5555, {N5104, N5260});
nand_n #(2, 0, 0) NAND_158 (N5562, {N5261, N5107});
nand_n #(2, 0, 0) NAND_159 (N5573, {N5262, N5109});
nand_n #(2, 0, 0) NAND_160 (N5579, {N5263, N5111});
nand_n #(2, 0, 0) NAND_161 (N5595, {N5274, N5114});
nand_n #(2, 0, 0) NAND_162 (N5606, {N5275, N5116});
nand_n #(2, 0, 0) NAND_163 (N5616, {N5180_0, N2715});
notg #(0, 0) NOT_329 (N5617, N5180_1);
notg #(0, 0) NOT_330 (N5618, N5183_0);
notg #(0, 0) NOT_331 (N5619, N5186_0);
notg #(0, 0) NOT_332 (N5620, N5189_0);
notg #(0, 0) NOT_333 (N5621, N5192_0);
notg #(0, 0) NOT_334 (N5622, N5195_0);
nand_n #(2, 0, 0) NAND_164 (N5624, {N5121, N5282});
nand_n #(2, 0, 0) NAND_165 (N5634, {N5123, N5283});
nand_n #(2, 0, 0) NAND_166 (N5655, {N5126, N5298});
nand_n #(2, 0, 0) NAND_167 (N5671, {N5128, N5299});
nand_n #(2, 0, 0) NAND_168 (N5684, {N5130, N5300});
notg #(0, 0) NOT_335 (N5690, N5202_0);
notg #(0, 0) NOT_336 (N5691, N5211_0);
nand_n #(2, 0, 0) NAND_169 (N5692, {N5303, N5304});
nand_n #(2, 0, 0) NAND_170 (N5696, {N5137, N5305});
nand_n #(2, 0, 0) NAND_171 (N5700, {N5306, N5140});
nand_n #(2, 0, 0) NAND_172 (N5703, {N5307, N5308});
nand_n #(2, 0, 0) NAND_173 (N5707, {N5309, N5310});
nand_n #(2, 0, 0) NAND_174 (N5711, {N5145, N5311});
and_n #(2, 0, 0) AND_416 (N5726, {N5166_0, N4512_1});
notg #(0, 0) NOT_337 (N5727, N5173_0);
notg #(0, 0) NOT_338 (N5728, N5177_0);
notg #(0, 0) NOT_339 (N5730, N5199_0);
notg #(0, 0) NOT_340 (N5731, N5205_0);
notg #(0, 0) NOT_341 (N5732, N5208_0);
notg #(0, 0) NOT_342 (N5733, N5214_0);
notg #(0, 0) NOT_343 (N5734, N5217_0);
notg #(0, 0) NOT_344 (N5735, N5220_0);
nand_n #(2, 0, 0) NAND_175 (N5736, {N5365, N5366});
nand_n #(2, 0, 0) NAND_176 (N5739, {N5363, N5364});
nand_n #(2, 0, 0) NAND_177 (N5742, {N5369, N5370});
nand_n #(2, 0, 0) NAND_178 (N5745, {N5367, N5368});
notg #(0, 0) NOT_345 (N5755, N5236_0);
nand_n #(2, 0, 0) NAND_179 (N5756, {N5332, N5331});
and_n #(2, 0, 0) AND_417 (N5954, {N5264_0, N4396_0});
nand_n #(2, 0, 0) NAND_180 (N5955, {N1899_1, N5617});
notg #(0, 0) NOT_346 (N5956, N5346_0);
and_n #(2, 0, 0) AND_418 (N6005, {N5284_0, N4456_0});
and_n #(2, 0, 0) AND_419 (N6006, {N5284_1, N4456_1});
notg #(0, 0) NOT_347 (N6023, N5371_0);
nand_n #(2, 0, 0) NAND_181 (N6024, {N5371_1, N5312});
notg #(0, 0) NOT_348 (N6025, N5315_0);
notg #(0, 0) NOT_349 (N6028, N5324_0);
bufg #(0, 0) BUF_255 (N6031, N5319_0);
bufg #(0, 0) BUF_256 (N6034, N5319_1);
bufg #(0, 0) BUF_257 (N6037, N5328_0);
bufg #(0, 0) BUF_258 (N6040, N5328_1);
notg #(0, 0) NOT_350 (N6044, N5385_0);
or_n #(2, 0, 0) OR_94 (N6045, {N5166_1, N5726});
bufg #(0, 0) BUF_259 (N6048, N5264_1);
bufg #(0, 0) BUF_260 (N6051, N5284_2);
bufg #(0, 0) BUF_261 (N6054, N5284_3);
notg #(0, 0) NOT_351 (N6065, N5374_0);
nand_n #(2, 0, 0) NAND_182 (N6066, {N5374_1, N5054});
notg #(0, 0) NOT_352 (N6067, N5377_0);
notg #(0, 0) NOT_353 (N6068, N5382_0);
nand_n #(2, 0, 0) NAND_183 (N6069, {N5382_1, N5755});
and_n #(2, 0, 0) AND_420 (N6071, {N5470_0, N4316_0});
and_n #(3, 0, 0) AND_421 (N6072, {N5477_0, N5470_1, N4320_0});
and_n #(4, 0, 0) AND_422 (N6073, {N5488_0, N5470_2, N4325_1, N5477_1});
and_n #(4, 0, 0) AND_423 (N6074, {N5562_0, N4357_4, N4385_1, N4364_5});
and_n #(2, 0, 0) AND_424 (N6075, {N5389_0, N4280_0});
and_n #(3, 0, 0) AND_425 (N6076, {N5396_0, N5389_1, N4284_0});
and_n #(4, 0, 0) AND_426 (N6077, {N5407_0, N5389_2, N4290_1, N5396_1});
and_n #(4, 0, 0) AND_427 (N6078, {N5624_0, N4418_4, N4445_1, N4425_5});
notg #(0, 0) NOT_354 (N6079, N5418_0);
and_n #(4, 0, 0) AND_428 (N6080, {N5396_2, N5418_1, N5407_1, N5389_3});
and_n #(2, 0, 0) AND_429 (N6083, {N5396_3, N4284_1});
and_n #(3, 0, 0) AND_430 (N6084, {N5407_2, N4290_2, N5396_4});
and_n #(3, 0, 0) AND_431 (N6085, {N5418_2, N5407_3, N5396_5});
and_n #(2, 0, 0) AND_432 (N6086, {N5396_6, N4284_2});
and_n #(3, 0, 0) AND_433 (N6087, {N4290_3, N5407_4, N5396_7});
and_n #(2, 0, 0) AND_434 (N6088, {N5407_5, N4290_4});
and_n #(2, 0, 0) AND_435 (N6089, {N5418_3, N5407_6});
and_n #(2, 0, 0) AND_436 (N6090, {N5407_7, N4290_5});
and_n #(5, 0, 0) AND_437 (N6091, {N5431_0, N5462_0, N5441_0, N5424_0, N5452_0});
and_n #(2, 0, 0) AND_438 (N6094, {N5424_1, N4298_0});
and_n #(3, 0, 0) AND_439 (N6095, {N5431_1, N5424_2, N4301_0});
and_n #(4, 0, 0) AND_440 (N6096, {N5441_1, N5424_3, N4305_0, N5431_2});
and_n #(5, 0, 0) AND_441 (N6097, {N5452_1, N5441_2, N5424_4, N4310_0, N5431_3});
and_n #(2, 0, 0) AND_442 (N6098, {N5431_4, N4301_1});
and_n #(3, 0, 0) AND_443 (N6099, {N5441_3, N4305_1, N5431_5});
and_n #(4, 0, 0) AND_444 (N6100, {N5452_2, N5441_4, N4310_1, N5431_6});
and_n #(5, 0, 0) AND_445 (N6101, {N4_1, N5462_1, N5441_5, N5452_3, N5431_7});
and_n #(2, 0, 0) AND_446 (N6102, {N4305_2, N5441_6});
and_n #(3, 0, 0) AND_447 (N6103, {N5452_4, N5441_7, N4310_2});
and_n #(4, 0, 0) AND_448 (N6104, {N4_2, N5462_2, N5441_8, N5452_5});
and_n #(2, 0, 0) AND_449 (N6105, {N5452_6, N4310_3});
and_n #(3, 0, 0) AND_450 (N6106, {N4_3, N5462_3, N5452_7});
and_n #(2, 0, 0) AND_451 (N6107, {N4_4, N5462_4});
and_n #(4, 0, 0) AND_452 (N6108, {N5549_0, N5488_1, N5477_2, N5470_3});
and_n #(2, 0, 0) AND_453 (N6111, {N5477_3, N4320_1});
and_n #(3, 0, 0) AND_454 (N6112, {N5488_2, N4325_2, N5477_4});
and_n #(3, 0, 0) AND_455 (N6113, {N5549_1, N5488_3, N5477_5});
and_n #(2, 0, 0) AND_456 (N6114, {N5477_6, N4320_2});
and_n #(3, 0, 0) AND_457 (N6115, {N5488_4, N4325_3, N5477_7});
and_n #(2, 0, 0) AND_458 (N6116, {N5488_5, N4325_4});
and_n #(5, 0, 0) AND_459 (N6117, {N5555_0, N5536_0, N5520_0, N5506_0, N5498_0});
and_n #(2, 0, 0) AND_460 (N6120, {N5498_1, N4332_0});
and_n #(3, 0, 0) AND_461 (N6121, {N5506_1, N5498_2, N4336_0});
and_n #(4, 0, 0) AND_462 (N6122, {N5520_1, N5498_3, N4342_0, N5506_2});
and_n #(5, 0, 0) AND_463 (N6123, {N5536_1, N5520_2, N5498_4, N4349_1, N5506_3});
and_n #(2, 0, 0) AND_464 (N6124, {N5506_4, N4336_1});
and_n #(3, 0, 0) AND_465 (N6125, {N5520_3, N4342_1, N5506_5});
and_n #(4, 0, 0) AND_466 (N6126, {N5536_2, N5520_4, N4349_2, N5506_6});
and_n #(4, 0, 0) AND_467 (N6127, {N5555_1, N5520_5, N5506_7, N5536_3});
and_n #(2, 0, 0) AND_468 (N6128, {N5506_8, N4336_2});
and_n #(3, 0, 0) AND_469 (N6129, {N5520_6, N4342_2, N5506_9});
and_n #(4, 0, 0) AND_470 (N6130, {N5536_4, N5520_7, N4349_3, N5506_10});
and_n #(2, 0, 0) AND_471 (N6131, {N5520_8, N4342_3});
and_n #(3, 0, 0) AND_472 (N6132, {N5536_5, N5520_9, N4349_4});
and_n #(3, 0, 0) AND_473 (N6133, {N5555_2, N5520_10, N5536_6});
and_n #(2, 0, 0) AND_474 (N6134, {N5520_11, N4342_4});
and_n #(3, 0, 0) AND_475 (N6135, {N5536_7, N5520_12, N4349_5});
and_n #(2, 0, 0) AND_476 (N6136, {N5536_8, N4349_6});
and_n #(2, 0, 0) AND_477 (N6137, {N5549_2, N5488_6});
and_n #(2, 0, 0) AND_478 (N6138, {N5555_3, N5536_9});
notg #(0, 0) NOT_355 (N6139, N5573_0);
and_n #(4, 0, 0) AND_479 (N6140, {N4364_6, N5573_1, N5562_1, N4357_5});
and_n #(3, 0, 0) AND_480 (N6143, {N5562_2, N4385_2, N4364_7});
and_n #(3, 0, 0) AND_481 (N6144, {N5573_2, N5562_3, N4364_8});
and_n #(3, 0, 0) AND_482 (N6145, {N4385_3, N5562_4, N4364_9});
and_n #(2, 0, 0) AND_483 (N6146, {N5562_5, N4385_4});
and_n #(2, 0, 0) AND_484 (N6147, {N5573_3, N5562_6});
and_n #(2, 0, 0) AND_485 (N6148, {N5562_7, N4385_5});
and_n #(5, 0, 0) AND_486 (N6149, {N5264_2, N4405_2, N5595_0, N5579_0, N5606_0});
and_n #(2, 0, 0) AND_487 (N6152, {N5579_1, N4067_0});
and_n #(3, 0, 0) AND_488 (N6153, {N5264_3, N5579_2, N4396_1});
and_n #(4, 0, 0) AND_489 (N6154, {N5595_1, N5579_3, N4400_0, N5264_4});
and_n #(5, 0, 0) AND_490 (N6155, {N5606_1, N5595_2, N5579_4, N4412_1, N5264_5});
and_n #(3, 0, 0) AND_491 (N6156, {N5595_3, N4400_1, N5264_6});
and_n #(4, 0, 0) AND_492 (N6157, {N5606_2, N5595_4, N4412_2, N5264_7});
and_n #(5, 0, 0) AND_493 (N6158, {N54_2, N4405_3, N5595_5, N5606_3, N5264_8});
and_n #(2, 0, 0) AND_494 (N6159, {N4400_2, N5595_6});
and_n #(3, 0, 0) AND_495 (N6160, {N5606_4, N5595_7, N4412_3});
and_n #(4, 0, 0) AND_496 (N6161, {N54_3, N4405_4, N5595_8, N5606_5});
and_n #(2, 0, 0) AND_497 (N6162, {N5606_6, N4412_4});
and_n #(3, 0, 0) AND_498 (N6163, {N54_4, N4405_5, N5606_7});
nand_n #(2, 0, 0) NAND_184 (N6164, {N5616, N5955});
and_n #(4, 0, 0) AND_499 (N6168, {N5684_0, N5624_1, N4425_6, N4418_5});
and_n #(3, 0, 0) AND_500 (N6171, {N5624_2, N4445_2, N4425_7});
and_n #(3, 0, 0) AND_501 (N6172, {N5684_1, N5624_3, N4425_8});
and_n #(3, 0, 0) AND_502 (N6173, {N5624_4, N4445_3, N4425_9});
and_n #(2, 0, 0) AND_503 (N6174, {N5624_5, N4445_4});
and_n #(5, 0, 0) AND_504 (N6175, {N4477_2, N5671_0, N5655_0, N5284_4, N5634_0});
and_n #(2, 0, 0) AND_505 (N6178, {N5634_1, N4080_0});
and_n #(3, 0, 0) AND_506 (N6179, {N5284_5, N5634_2, N4456_2});
and_n #(4, 0, 0) AND_507 (N6180, {N5655_1, N5634_3, N4462_0, N5284_6});
and_n #(5, 0, 0) AND_508 (N6181, {N5671_1, N5655_2, N5634_4, N4469_1, N5284_7});
and_n #(3, 0, 0) AND_509 (N6182, {N5655_3, N4462_1, N5284_8});
and_n #(4, 0, 0) AND_510 (N6183, {N5671_2, N5655_4, N4469_2, N5284_9});
and_n #(4, 0, 0) AND_511 (N6184, {N4477_3, N5655_5, N5284_10, N5671_3});
and_n #(3, 0, 0) AND_512 (N6185, {N5655_6, N4462_2, N5284_11});
and_n #(4, 0, 0) AND_513 (N6186, {N5671_4, N5655_7, N4469_3, N5284_12});
and_n #(2, 0, 0) AND_514 (N6187, {N5655_8, N4462_3});
and_n #(3, 0, 0) AND_515 (N6188, {N5671_5, N5655_9, N4469_4});
and_n #(3, 0, 0) AND_516 (N6189, {N4477_4, N5655_10, N5671_6});
and_n #(2, 0, 0) AND_517 (N6190, {N5655_11, N4462_4});
and_n #(3, 0, 0) AND_518 (N6191, {N5671_7, N5655_12, N4469_5});
and_n #(2, 0, 0) AND_519 (N6192, {N5671_8, N4469_6});
and_n #(2, 0, 0) AND_520 (N6193, {N5684_2, N5624_6});
and_n #(2, 0, 0) AND_521 (N6194, {N4477_5, N5671_9});
notg #(0, 0) NOT_356 (N6197, N5692_0);
notg #(0, 0) NOT_357 (N6200, N5696_0);
notg #(0, 0) NOT_358 (N6203, N5703_0);
notg #(0, 0) NOT_359 (N6206, N5707_0);
bufg #(0, 0) BUF_262 (N6209, N5700_0);
bufg #(0, 0) BUF_263 (N6212, N5700_1);
bufg #(0, 0) BUF_264 (N6215, N5711_0);
bufg #(0, 0) BUF_265 (N6218, N5711_1);
nand_n #(2, 0, 0) NAND_185 (N6221, {N5049_1, N6023});
notg #(0, 0) NOT_360 (N6234, N5756_0);
nand_n #(2, 0, 0) NAND_186 (N6235, {N5756_1, N6044});
bufg #(0, 0) BUF_266 (N6238, N5462_5);
bufg #(0, 0) BUF_267 (N6241, N5389_4);
bufg #(0, 0) BUF_268 (N6244, N5389_5);
bufg #(0, 0) BUF_269 (N6247, N5396_8);
bufg #(0, 0) BUF_270 (N6250, N5396_9);
bufg #(0, 0) BUF_271 (N6253, N5407_8);
bufg #(0, 0) BUF_272 (N6256, N5407_9);
bufg #(0, 0) BUF_273 (N6259, N5424_5);
bufg #(0, 0) BUF_274 (N6262, N5431_8);
bufg #(0, 0) BUF_275 (N6265, N5441_9);
bufg #(0, 0) BUF_276 (N6268, N5452_8);
bufg #(0, 0) BUF_277 (N6271, N5549_3);
bufg #(0, 0) BUF_278 (N6274, N5488_7);
bufg #(0, 0) BUF_279 (N6277, N5470_4);
bufg #(0, 0) BUF_280 (N6280, N5477_8);
bufg #(0, 0) BUF_281 (N6283, N5549_4);
bufg #(0, 0) BUF_282 (N6286, N5488_8);
bufg #(0, 0) BUF_283 (N6289, N5470_5);
bufg #(0, 0) BUF_284 (N6292, N5477_9);
bufg #(0, 0) BUF_285 (N6295, N5555_4);
bufg #(0, 0) BUF_286 (N6298, N5536_10);
bufg #(0, 0) BUF_287 (N6301, N5498_5);
bufg #(0, 0) BUF_288 (N6304, N5520_13);
bufg #(0, 0) BUF_289 (N6307, N5506_11);
bufg #(0, 0) BUF_290 (N6310, N5506_12);
bufg #(0, 0) BUF_291 (N6313, N5555_5);
bufg #(0, 0) BUF_292 (N6316, N5536_11);
bufg #(0, 0) BUF_293 (N6319, N5498_6);
bufg #(0, 0) BUF_294 (N6322, N5520_14);
bufg #(0, 0) BUF_295 (N6325, N5562_8);
bufg #(0, 0) BUF_296 (N6328, N5562_9);
bufg #(0, 0) BUF_297 (N6331, N5579_5);
bufg #(0, 0) BUF_298 (N6335, N5595_9);
bufg #(0, 0) BUF_299 (N6338, N5606_8);
bufg #(0, 0) BUF_300 (N6341, N5684_3);
bufg #(0, 0) BUF_301 (N6344, N5624_7);
bufg #(0, 0) BUF_302 (N6347, N5684_4);
bufg #(0, 0) BUF_303 (N6350, N5624_8);
bufg #(0, 0) BUF_304 (N6353, N5671_10);
bufg #(0, 0) BUF_305 (N6356, N5634_5);
bufg #(0, 0) BUF_306 (N6359, N5655_13);
bufg #(0, 0) BUF_307 (N6364, N5671_11);
bufg #(0, 0) BUF_308 (N6367, N5634_6);
bufg #(0, 0) BUF_309 (N6370, N5655_14);
notg #(0, 0) NOT_361 (N6373, N5736_0);
notg #(0, 0) NOT_362 (N6374, N5739_0);
notg #(0, 0) NOT_363 (N6375, N5742_0);
notg #(0, 0) NOT_364 (N6376, N5745_0);
nand_n #(2, 0, 0) NAND_187 (N6377, {N4243_1, N6065});
nand_n #(2, 0, 0) NAND_188 (N6378, {N5236_1, N6068});
or_n #(4, 0, 0) OR_95 (N6382, {N4268, N6071, N6072, N6073});
or_n #(4, 0, 0) OR_96 (N6386, {N3968_4, N5065, N5066, N6074});
or_n #(4, 0, 0) OR_97 (N6388, {N4271, N6075, N6076, N6077});
or_n #(4, 0, 0) OR_98 (N6392, {N3968_5, N5067, N5068, N6078});
or_n #(5, 0, 0) OR_99 (N6397, {N4297, N6094, N6095, N6096, N6097});
or_n #(2, 0, 0) OR_100 (N6411, {N4320_3, N6116});
or_n #(5, 0, 0) OR_101 (N6415, {N4331, N6120, N6121, N6122, N6123});
or_n #(2, 0, 0) OR_102 (N6419, {N4342_5, N6136});
or_n #(5, 0, 0) OR_103 (N6427, {N4392, N6152, N6153, N6154, N6155});
notg #(0, 0) NOT_365 (N6434, N6048_0);
or_n #(2, 0, 0) OR_104 (N6437, {N4440_3, N6174});
or_n #(5, 0, 0) OR_105 (N6441, {N4451, N6178, N6179, N6180, N6181});
or_n #(2, 0, 0) OR_106 (N6445, {N4462_5, N6192});
notg #(0, 0) NOT_366 (N6448, N6051_0);
notg #(0, 0) NOT_367 (N6449, N6054_0);
nand_n #(2, 0, 0) NAND_189 (N6466, {N6221, N6024});
notg #(0, 0) NOT_368 (N6469, N6031_0);
notg #(0, 0) NOT_369 (N6470, N6034_0);
notg #(0, 0) NOT_370 (N6471, N6037_0);
notg #(0, 0) NOT_371 (N6472, N6040_0);
and_n #(3, 0, 0) AND_522 (N6473, {N5315_1, N4524_1, N6031_1});
and_n #(3, 0, 0) AND_523 (N6474, {N6025_0, N5150_0, N6034_1});
and_n #(3, 0, 0) AND_524 (N6475, {N5324_1, N4532_1, N6037_1});
and_n #(3, 0, 0) AND_525 (N6476, {N6028_0, N5157_0, N6040_1});
nand_n #(2, 0, 0) NAND_190 (N6477, {N5385_1, N6234});
nand_n #(2, 0, 0) NAND_191 (N6478, {N6045_0, N132_0});
or_n #(4, 0, 0) OR_107 (N6482, {N4280_1, N6083, N6084, N6085});
nor_n #(3, 0, 0) NOR_10 (N6486, {N4280_2, N6086, N6087});
or_n #(3, 0, 0) OR_108 (N6490, {N4284_3, N6088, N6089});
nor_n #(2, 0, 0) NOR_11 (N6494, {N4284_4, N6090});
or_n #(5, 0, 0) OR_109 (N6500, {N4298_1, N6098, N6099, N6100, N6101});
or_n #(4, 0, 0) OR_110 (N6504, {N4301_2, N6102, N6103, N6104});
or_n #(3, 0, 0) OR_111 (N6508, {N4305_3, N6105, N6106});
or_n #(2, 0, 0) OR_112 (N6512, {N4310_4, N6107});
or_n #(4, 0, 0) OR_113 (N6516, {N4316_1, N6111, N6112, N6113});
nor_n #(3, 0, 0) NOR_12 (N6526, {N4316_2, N6114, N6115});
or_n #(4, 0, 0) OR_114 (N6536, {N4336_3, N6131, N6132, N6133});
or_n #(5, 0, 0) OR_115 (N6539, {N4332_1, N6124, N6125, N6126, N6127});
nor_n #(3, 0, 0) NOR_13 (N6553, {N4336_4, N6134, N6135});
nor_n #(4, 0, 0) NOR_14 (N6556, {N4332_2, N6128, N6129, N6130});
or_n #(4, 0, 0) OR_116 (N6566, {N4375_1, N5117, N6143, N6144});
nor_n #(3, 0, 0) NOR_15 (N6569, {N4375_2, N5118, N6145});
or_n #(3, 0, 0) OR_117 (N6572, {N4379_3, N6146, N6147});
nor_n #(2, 0, 0) NOR_16 (N6575, {N4379_4, N6148});
or_n #(5, 0, 0) OR_118 (N6580, {N4067_1, N5954, N6156, N6157, N6158});
or_n #(4, 0, 0) OR_119 (N6584, {N4396_2, N6159, N6160, N6161});
or_n #(3, 0, 0) OR_120 (N6587, {N4400_3, N6162, N6163});
or_n #(4, 0, 0) OR_121 (N6592, {N4436_1, N5132, N6171, N6172});
nor_n #(3, 0, 0) NOR_17 (N6599, {N4436_2, N5133, N6173});
or_n #(4, 0, 0) OR_122 (N6606, {N4456_3, N6187, N6188, N6189});
or_n #(5, 0, 0) OR_123 (N6609, {N4080_1, N6005, N6182, N6183, N6184});
nor_n #(3, 0, 0) NOR_18 (N6619, {N4456_4, N6190, N6191});
nor_n #(4, 0, 0) NOR_19 (N6622, {N4080_2, N6006, N6185, N6186});
nand_n #(2, 0, 0) NAND_192 (N6630, {N5739_1, N6373});
nand_n #(2, 0, 0) NAND_193 (N6631, {N5736_1, N6374});
nand_n #(2, 0, 0) NAND_194 (N6632, {N5745_1, N6375});
nand_n #(2, 0, 0) NAND_195 (N6633, {N5742_1, N6376});
nand_n #(2, 0, 0) NAND_196 (N6634, {N6377, N6066});
nand_n #(2, 0, 0) NAND_197 (N6637, {N6069, N6378});
notg #(0, 0) NOT_372 (N6640, N6164_0);
and_n #(2, 0, 0) AND_526 (N6641, {N6108_0, N6117_0});
and_n #(2, 0, 0) AND_527 (N6643, {N6140_0, N6149_0});
and_n #(2, 0, 0) AND_528 (N6646, {N6168_0, N6175_0});
and_n #(2, 0, 0) AND_529 (N6648, {N6080_0, N6091_0});
nand_n #(2, 0, 0) NAND_198 (N6650, {N6238_0, N2637});
notg #(0, 0) NOT_373 (N6651, N6238_1);
notg #(0, 0) NOT_374 (N6653, N6241_0);
notg #(0, 0) NOT_375 (N6655, N6244_0);
notg #(0, 0) NOT_376 (N6657, N6247_0);
notg #(0, 0) NOT_377 (N6659, N6250_0);
nand_n #(2, 0, 0) NAND_199 (N6660, {N6253_0, N5087});
notg #(0, 0) NOT_378 (N6661, N6253_1);
nand_n #(2, 0, 0) NAND_200 (N6662, {N6256_0, N5469});
notg #(0, 0) NOT_379 (N6663, N6256_1);
and_n #(2, 0, 0) AND_530 (N6664, {N6091_1, N4_5});
notg #(0, 0) NOT_380 (N6666, N6259_0);
notg #(0, 0) NOT_381 (N6668, N6262_0);
notg #(0, 0) NOT_382 (N6670, N6265_0);
notg #(0, 0) NOT_383 (N6672, N6268_0);
notg #(0, 0) NOT_384 (N6675, N6117_1);
notg #(0, 0) NOT_385 (N6680, N6280_0);
notg #(0, 0) NOT_386 (N6681, N6292_0);
notg #(0, 0) NOT_387 (N6682, N6307_0);
notg #(0, 0) NOT_388 (N6683, N6310_0);
nand_n #(2, 0, 0) NAND_201 (N6689, {N6325_0, N5120});
notg #(0, 0) NOT_389 (N6690, N6325_1);
nand_n #(2, 0, 0) NAND_202 (N6691, {N6328_0, N5622});
notg #(0, 0) NOT_390 (N6692, N6328_1);
and_n #(2, 0, 0) AND_531 (N6693, {N6149_1, N54_5});
notg #(0, 0) NOT_391 (N6695, N6331_0);
notg #(0, 0) NOT_392 (N6698, N6335_0);
nand_n #(2, 0, 0) NAND_203 (N6699, {N6338_0, N5956});
notg #(0, 0) NOT_393 (N6700, N6338_1);
notg #(0, 0) NOT_394 (N6703, N6175_1);
notg #(0, 0) NOT_395 (N6708, N6209_0);
notg #(0, 0) NOT_396 (N6709, N6212_0);
notg #(0, 0) NOT_397 (N6710, N6215_0);
notg #(0, 0) NOT_398 (N6711, N6218_0);
and_n #(3, 0, 0) AND_532 (N6712, {N5696_1, N5692_1, N6209_1});
and_n #(3, 0, 0) AND_533 (N6713, {N6200_0, N6197_0, N6212_1});
and_n #(3, 0, 0) AND_534 (N6714, {N5707_1, N5703_1, N6215_1});
and_n #(3, 0, 0) AND_535 (N6715, {N6206_0, N6203_0, N6218_1});
bufg #(0, 0) BUF_310 (N6716, N6466_0);
and_n #(3, 0, 0) AND_536 (N6718, {N6164_1, N1777_2, N3130_4});
and_n #(3, 0, 0) AND_537 (N6719, {N5150_1, N5315_2, N6469});
and_n #(3, 0, 0) AND_538 (N6720, {N4524_2, N6025_1, N6470});
and_n #(3, 0, 0) AND_539 (N6721, {N5157_1, N5324_2, N6471});
and_n #(3, 0, 0) AND_540 (N6722, {N4532_2, N6028_1, N6472});
nand_n #(2, 0, 0) NAND_204 (N6724, {N6477, N6235});
notg #(0, 0) NOT_399 (N6739, N6271_0);
notg #(0, 0) NOT_400 (N6740, N6274_0);
notg #(0, 0) NOT_401 (N6741, N6277_0);
notg #(0, 0) NOT_402 (N6744, N6283_0);
notg #(0, 0) NOT_403 (N6745, N6286_0);
notg #(0, 0) NOT_404 (N6746, N6289_0);
notg #(0, 0) NOT_405 (N6751, N6295_0);
notg #(0, 0) NOT_406 (N6752, N6298_0);
notg #(0, 0) NOT_407 (N6753, N6301_0);
notg #(0, 0) NOT_408 (N6754, N6304_0);
notg #(0, 0) NOT_409 (N6755, N6322_0);
notg #(0, 0) NOT_410 (N6760, N6313_0);
notg #(0, 0) NOT_411 (N6761, N6316_0);
notg #(0, 0) NOT_412 (N6762, N6319_0);
notg #(0, 0) NOT_413 (N6772, N6341_0);
notg #(0, 0) NOT_414 (N6773, N6344_0);
notg #(0, 0) NOT_415 (N6776, N6347_0);
notg #(0, 0) NOT_416 (N6777, N6350_0);
notg #(0, 0) NOT_417 (N6782, N6353_0);
notg #(0, 0) NOT_418 (N6783, N6356_0);
notg #(0, 0) NOT_419 (N6784, N6359_0);
notg #(0, 0) NOT_420 (N6785, N6370_0);
notg #(0, 0) NOT_421 (N6790, N6364_0);
notg #(0, 0) NOT_422 (N6791, N6367_0);
nand_n #(2, 0, 0) NAND_205 (N6792, {N6630, N6631});
nand_n #(2, 0, 0) NAND_206 (N6795, {N6632, N6633});
and_n #(2, 0, 0) AND_541 (N6801, {N6108_1, N6415_0});
and_n #(2, 0, 0) AND_542 (N6802, {N6427_0, N6140_1});
and_n #(2, 0, 0) AND_543 (N6803, {N6397_0, N6080_1});
and_n #(2, 0, 0) AND_544 (N6804, {N6168_1, N6441_0});
notg #(0, 0) NOT_423 (N6805, N6466_1);
nand_n #(2, 0, 0) NAND_207 (N6806, {N1851_1, N6651});
notg #(0, 0) NOT_424 (N6807, N6482_0);
nand_n #(2, 0, 0) NAND_208 (N6808, {N6482_1, N6653});
notg #(0, 0) NOT_425 (N6809, N6486_0);
nand_n #(2, 0, 0) NAND_209 (N6810, {N6486_1, N6655});
notg #(0, 0) NOT_426 (N6811, N6490_0);
nand_n #(2, 0, 0) NAND_210 (N6812, {N6490_1, N6657});
notg #(0, 0) NOT_427 (N6813, N6494_0);
nand_n #(2, 0, 0) NAND_211 (N6814, {N6494_1, N6659});
nand_n #(2, 0, 0) NAND_212 (N6815, {N4575_1, N6661});
nand_n #(2, 0, 0) NAND_213 (N6816, {N5169_1, N6663});
or_n #(2, 0, 0) OR_124 (N6817, {N6397_1, N6664});
notg #(0, 0) NOT_428 (N6823, N6500_0);
nand_n #(2, 0, 0) NAND_214 (N6824, {N6500_1, N6666});
notg #(0, 0) NOT_429 (N6825, N6504_0);
nand_n #(2, 0, 0) NAND_215 (N6826, {N6504_1, N6668});
notg #(0, 0) NOT_430 (N6827, N6508_0);
nand_n #(2, 0, 0) NAND_216 (N6828, {N6508_1, N6670});
notg #(0, 0) NOT_431 (N6829, N6512_0);
nand_n #(2, 0, 0) NAND_217 (N6830, {N6512_1, N6672});
notg #(0, 0) NOT_432 (N6831, N6415_1);
notg #(0, 0) NOT_433 (N6834, N6566_0);
nand_n #(2, 0, 0) NAND_218 (N6835, {N6566_1, N5618});
notg #(0, 0) NOT_434 (N6836, N6569_0);
nand_n #(2, 0, 0) NAND_219 (N6837, {N6569_1, N5619});
notg #(0, 0) NOT_435 (N6838, N6572_0);
nand_n #(2, 0, 0) NAND_220 (N6839, {N6572_1, N5620});
notg #(0, 0) NOT_436 (N6840, N6575_0);
nand_n #(2, 0, 0) NAND_221 (N6841, {N6575_1, N5621});
nand_n #(2, 0, 0) NAND_222 (N6842, {N4627_1, N6690});
nand_n #(2, 0, 0) NAND_223 (N6843, {N5195_1, N6692});
or_n #(2, 0, 0) OR_125 (N6844, {N6427_1, N6693});
notg #(0, 0) NOT_437 (N6850, N6580_0);
nand_n #(2, 0, 0) NAND_224 (N6851, {N6580_1, N6695});
notg #(0, 0) NOT_438 (N6852, N6584_0);
nand_n #(2, 0, 0) NAND_225 (N6853, {N6584_1, N6434});
notg #(0, 0) NOT_439 (N6854, N6587_0);
nand_n #(2, 0, 0) NAND_226 (N6855, {N6587_1, N6698});
nand_n #(2, 0, 0) NAND_227 (N6856, {N5346_1, N6700});
notg #(0, 0) NOT_440 (N6857, N6441_1);
and_n #(3, 0, 0) AND_545 (N6860, {N6197_1, N5696_2, N6708});
and_n #(3, 0, 0) AND_546 (N6861, {N5692_2, N6200_1, N6709});
and_n #(3, 0, 0) AND_547 (N6862, {N6203_1, N5707_2, N6710});
and_n #(3, 0, 0) AND_548 (N6863, {N5703_2, N6206_1, N6711});
or_n #(3, 0, 0) OR_126 (N6866, {N4197, N6718, N3785});
nor_n #(2, 0, 0) NOR_20 (N6872, {N6719, N6473});
nor_n #(2, 0, 0) NOR_21 (N6873, {N6720, N6474});
nor_n #(2, 0, 0) NOR_22 (N6874, {N6721, N6475});
nor_n #(2, 0, 0) NOR_23 (N6875, {N6722, N6476});
notg #(0, 0) NOT_441 (N6876, N6637_0);
bufg #(0, 0) BUF_311 (N6877, N6724_0);
and_n #(2, 0, 0) AND_549 (N6879, {N6045_1, N6478_0});
and_n #(2, 0, 0) AND_550 (N6880, {N6478_1, N132_1});
or_n #(2, 0, 0) OR_127 (N6881, {N6411_0, N6137});
notg #(0, 0) NOT_442 (N6884, N6516_0);
notg #(0, 0) NOT_443 (N6885, N6411_1);
notg #(0, 0) NOT_444 (N6888, N6526_0);
notg #(0, 0) NOT_445 (N6889, N6536_0);
nand_n #(2, 0, 0) NAND_228 (N6890, {N6536_1, N5176});
or_n #(2, 0, 0) OR_128 (N6891, {N6419_0, N6138});
notg #(0, 0) NOT_446 (N6894, N6539_0);
notg #(0, 0) NOT_447 (N6895, N6553_0);
nand_n #(2, 0, 0) NAND_229 (N6896, {N6553_1, N5728});
notg #(0, 0) NOT_448 (N6897, N6419_1);
notg #(0, 0) NOT_449 (N6900, N6556_0);
or_n #(2, 0, 0) OR_129 (N6901, {N6437_0, N6193});
notg #(0, 0) NOT_450 (N6904, N6592_0);
notg #(0, 0) NOT_451 (N6905, N6437_1);
notg #(0, 0) NOT_452 (N6908, N6599_0);
or_n #(2, 0, 0) OR_130 (N6909, {N6445_0, N6194});
notg #(0, 0) NOT_453 (N6912, N6606_0);
notg #(0, 0) NOT_454 (N6913, N6609_0);
notg #(0, 0) NOT_455 (N6914, N6619_0);
nand_n #(2, 0, 0) NAND_230 (N6915, {N6619_1, N5734});
notg #(0, 0) NOT_456 (N6916, N6445_1);
notg #(0, 0) NOT_457 (N6919, N6622_0);
notg #(0, 0) NOT_458 (N6922, N6634_0);
nand_n #(2, 0, 0) NAND_231 (N6923, {N6634_1, N6067});
or_n #(2, 0, 0) OR_131 (N6924, {N6382, N6801});
or_n #(2, 0, 0) OR_132 (N6925, {N6386, N6802});
or_n #(2, 0, 0) OR_133 (N6926, {N6388, N6803});
or_n #(2, 0, 0) OR_134 (N6927, {N6392, N6804});
notg #(0, 0) NOT_459 (N6930, N6724_1);
nand_n #(2, 0, 0) NAND_232 (N6932, {N6650, N6806});
nand_n #(2, 0, 0) NAND_233 (N6935, {N6241_1, N6807});
nand_n #(2, 0, 0) NAND_234 (N6936, {N6244_1, N6809});
nand_n #(2, 0, 0) NAND_235 (N6937, {N6247_1, N6811});
nand_n #(2, 0, 0) NAND_236 (N6938, {N6250_1, N6813});
nand_n #(2, 0, 0) NAND_237 (N6939, {N6660, N6815});
nand_n #(2, 0, 0) NAND_238 (N6940, {N6662, N6816});
nand_n #(2, 0, 0) NAND_239 (N6946, {N6259_1, N6823});
nand_n #(2, 0, 0) NAND_240 (N6947, {N6262_1, N6825});
nand_n #(2, 0, 0) NAND_241 (N6948, {N6265_1, N6827});
nand_n #(2, 0, 0) NAND_242 (N6949, {N6268_1, N6829});
nand_n #(2, 0, 0) NAND_243 (N6953, {N5183_1, N6834});
nand_n #(2, 0, 0) NAND_244 (N6954, {N5186_1, N6836});
nand_n #(2, 0, 0) NAND_245 (N6955, {N5189_1, N6838});
nand_n #(2, 0, 0) NAND_246 (N6956, {N5192_1, N6840});
nand_n #(2, 0, 0) NAND_247 (N6957, {N6689, N6842});
nand_n #(2, 0, 0) NAND_248 (N6958, {N6691, N6843});
nand_n #(2, 0, 0) NAND_249 (N6964, {N6331_1, N6850});
nand_n #(2, 0, 0) NAND_250 (N6965, {N6048_1, N6852});
nand_n #(2, 0, 0) NAND_251 (N6966, {N6335_1, N6854});
nand_n #(2, 0, 0) NAND_252 (N6967, {N6699, N6856});
nor_n #(2, 0, 0) NOR_24 (N6973, {N6860, N6712});
nor_n #(2, 0, 0) NOR_25 (N6974, {N6861, N6713});
nor_n #(2, 0, 0) NOR_26 (N6975, {N6862, N6714});
nor_n #(2, 0, 0) NOR_27 (N6976, {N6863, N6715});
notg #(0, 0) NOT_460 (N6977, N6792_0);
notg #(0, 0) NOT_461 (N6978, N6795_0);
or_n #(2, 0, 0) OR_135 (N6979, {N6879, N6880});
nand_n #(2, 0, 0) NAND_253 (N6987, {N4608_1, N6889});
nand_n #(2, 0, 0) NAND_254 (N6990, {N5177_1, N6895});
nand_n #(2, 0, 0) NAND_255 (N6999, {N5217_1, N6914});
nand_n #(2, 0, 0) NAND_256 (N7002, {N5377_1, N6922});
nand_n #(2, 0, 0) NAND_257 (N7003, {N6873, N6872});
nand_n #(2, 0, 0) NAND_258 (N7006, {N6875, N6874});
and_n #(3, 0, 0) AND_551 (N7011, {N6866_0, N2681_5, N2692_0});
and_n #(3, 0, 0) AND_552 (N7012, {N6866_1, N2756_5, N2767_0});
and_n #(3, 0, 0) AND_553 (N7013, {N6866_2, N2779_5, N2790_0});
notg #(0, 0) NOT_462 (N7015, N6866_3);
and_n #(3, 0, 0) AND_554 (N7016, {N6866_4, N2801_5, N2812_0});
nand_n #(2, 0, 0) NAND_259 (N7018, {N6935, N6808});
nand_n #(2, 0, 0) NAND_260 (N7019, {N6936, N6810});
nand_n #(2, 0, 0) NAND_261 (N7020, {N6937, N6812});
nand_n #(2, 0, 0) NAND_262 (N7021, {N6938, N6814});
notg #(0, 0) NOT_463 (N7022, N6939);
notg #(0, 0) NOT_464 (N7023, N6817_0);
nand_n #(2, 0, 0) NAND_263 (N7028, {N6946, N6824});
nand_n #(2, 0, 0) NAND_264 (N7031, {N6947, N6826});
nand_n #(2, 0, 0) NAND_265 (N7034, {N6948, N6828});
nand_n #(2, 0, 0) NAND_266 (N7037, {N6949, N6830});
and_n #(2, 0, 0) AND_555 (N7040, {N6817_1, N6079});
and_n #(2, 0, 0) AND_556 (N7041, {N6831_0, N6675});
nand_n #(2, 0, 0) NAND_267 (N7044, {N6953, N6835});
nand_n #(2, 0, 0) NAND_268 (N7045, {N6954, N6837});
nand_n #(2, 0, 0) NAND_269 (N7046, {N6955, N6839});
nand_n #(2, 0, 0) NAND_270 (N7047, {N6956, N6841});
notg #(0, 0) NOT_465 (N7048, N6957);
notg #(0, 0) NOT_466 (N7049, N6844_0);
nand_n #(2, 0, 0) NAND_271 (N7054, {N6964, N6851});
nand_n #(2, 0, 0) NAND_272 (N7057, {N6965, N6853});
nand_n #(2, 0, 0) NAND_273 (N7060, {N6966, N6855});
and_n #(2, 0, 0) AND_557 (N7064, {N6844_1, N6139});
and_n #(2, 0, 0) AND_558 (N7065, {N6857_0, N6703});
notg #(0, 0) NOT_467 (N7072, N6881_0);
nand_n #(2, 0, 0) NAND_274 (N7073, {N6881_1, N5172});
notg #(0, 0) NOT_468 (N7074, N6885_0);
nand_n #(2, 0, 0) NAND_275 (N7075, {N6885_1, N5727});
nand_n #(2, 0, 0) NAND_276 (N7076, {N6890, N6987});
notg #(0, 0) NOT_469 (N7079, N6891_0);
nand_n #(2, 0, 0) NAND_277 (N7080, {N6896, N6990});
notg #(0, 0) NOT_470 (N7083, N6897_0);
notg #(0, 0) NOT_471 (N7084, N6901_0);
nand_n #(2, 0, 0) NAND_278 (N7085, {N6901_1, N5198});
notg #(0, 0) NOT_472 (N7086, N6905_0);
nand_n #(2, 0, 0) NAND_279 (N7087, {N6905_1, N5731});
notg #(0, 0) NOT_473 (N7088, N6909_0);
nand_n #(2, 0, 0) NAND_280 (N7089, {N6909_1, N6912});
nand_n #(2, 0, 0) NAND_281 (N7090, {N6915, N6999});
notg #(0, 0) NOT_474 (N7093, N6916_0);
nand_n #(2, 0, 0) NAND_282 (N7094, {N6974, N6973});
nand_n #(2, 0, 0) NAND_283 (N7097, {N6976, N6975});
nand_n #(2, 0, 0) NAND_284 (N7101, {N7002, N6923});
notg #(0, 0) NOT_475 (N7105, N6932_0);
notg #(0, 0) NOT_476 (N7110, N6967_0);
and_n #(3, 0, 0) AND_559 (N7114, {N6979_0, N603_1, N1755_1});
notg #(0, 0) NOT_477 (N7115, N7019);
notg #(0, 0) NOT_478 (N7116, N7021);
and_n #(2, 0, 0) AND_560 (N7125, {N6817_2, N7018});
and_n #(2, 0, 0) AND_561 (N7126, {N6817_3, N7020});
and_n #(2, 0, 0) AND_562 (N7127, {N6817_4, N7022});
notg #(0, 0) NOT_479 (N7130, N7045);
notg #(0, 0) NOT_480 (N7131, N7047);
and_n #(2, 0, 0) AND_563 (N7139, {N6844_2, N7044});
and_n #(2, 0, 0) AND_564 (N7140, {N6844_3, N7046});
and_n #(2, 0, 0) AND_565 (N7141, {N6844_4, N7048});
and_n #(3, 0, 0) AND_566 (N7146, {N6932_1, N1761_2, N3108_4});
and_n #(3, 0, 0) AND_567 (N7147, {N6967_1, N1777_3, N3130_5});
notg #(0, 0) NOT_481 (N7149, N7003_0);
notg #(0, 0) NOT_482 (N7150, N7006_0);
nand_n #(2, 0, 0) NAND_285 (N7151, {N7006_1, N6876});
nand_n #(2, 0, 0) NAND_286 (N7152, {N4605_1, N7072});
nand_n #(2, 0, 0) NAND_287 (N7153, {N5173_1, N7074});
nand_n #(2, 0, 0) NAND_288 (N7158, {N4646_1, N7084});
nand_n #(2, 0, 0) NAND_289 (N7159, {N5205_1, N7086});
nand_n #(2, 0, 0) NAND_290 (N7160, {N6606_1, N7088});
notg #(0, 0) NOT_483 (N7166, N7037_0);
notg #(0, 0) NOT_484 (N7167, N7034_0);
notg #(0, 0) NOT_485 (N7168, N7031_0);
notg #(0, 0) NOT_486 (N7169, N7028_0);
notg #(0, 0) NOT_487 (N7170, N7060_0);
notg #(0, 0) NOT_488 (N7171, N7057_0);
notg #(0, 0) NOT_489 (N7172, N7054_0);
and_n #(2, 0, 0) AND_568 (N7173, {N7115, N7023_0});
and_n #(2, 0, 0) AND_569 (N7174, {N7116, N7023_1});
and_n #(2, 0, 0) AND_570 (N7175, {N6940, N7023_2});
and_n #(2, 0, 0) AND_571 (N7176, {N5418_4, N7023_3});
notg #(0, 0) NOT_490 (N7177, N7041_0);
and_n #(2, 0, 0) AND_572 (N7178, {N7130, N7049_0});
and_n #(2, 0, 0) AND_573 (N7179, {N7131, N7049_1});
and_n #(2, 0, 0) AND_574 (N7180, {N6958, N7049_2});
and_n #(2, 0, 0) AND_575 (N7181, {N5573_4, N7049_3});
notg #(0, 0) NOT_491 (N7182, N7065_0);
notg #(0, 0) NOT_492 (N7183, N7094_0);
nand_n #(2, 0, 0) NAND_291 (N7184, {N7094_1, N6977});
notg #(0, 0) NOT_493 (N7185, N7097_0);
nand_n #(2, 0, 0) NAND_292 (N7186, {N7097_1, N6978});
and_n #(3, 0, 0) AND_576 (N7187, {N7037_1, N1761_3, N3108_5});
and_n #(3, 0, 0) AND_577 (N7188, {N7034_1, N1761_4, N3108_6});
and_n #(3, 0, 0) AND_578 (N7189, {N7031_1, N1761_5, N3108_7});
or_n #(3, 0, 0) OR_136 (N7190, {N4956, N7146, N3781});
and_n #(3, 0, 0) AND_579 (N7196, {N7060_1, N1777_4, N3130_6});
and_n #(3, 0, 0) AND_580 (N7197, {N7057_1, N1777_5, N3130_7});
or_n #(3, 0, 0) OR_137 (N7198, {N4960, N7147, N3786});
nand_n #(2, 0, 0) NAND_293 (N7204, {N7101_0, N7149});
notg #(0, 0) NOT_494 (N7205, N7101_1);
nand_n #(2, 0, 0) NAND_294 (N7206, {N6637_1, N7150});
and_n #(3, 0, 0) AND_581 (N7207, {N7028_1, N1793_1, N3158_5});
and_n #(3, 0, 0) AND_582 (N7208, {N7054_1, N1807_1, N3180_5});
nand_n #(2, 0, 0) NAND_295 (N7209, {N7073, N7152});
nand_n #(2, 0, 0) NAND_296 (N7212, {N7075, N7153});
notg #(0, 0) NOT_495 (N7215, N7076_0);
nand_n #(2, 0, 0) NAND_297 (N7216, {N7076_1, N7079});
notg #(0, 0) NOT_496 (N7217, N7080_0);
nand_n #(2, 0, 0) NAND_298 (N7218, {N7080_1, N7083});
nand_n #(2, 0, 0) NAND_299 (N7219, {N7085, N7158});
nand_n #(2, 0, 0) NAND_300 (N7222, {N7087, N7159});
nand_n #(2, 0, 0) NAND_301 (N7225, {N7089, N7160});
notg #(0, 0) NOT_497 (N7228, N7090_0);
nand_n #(2, 0, 0) NAND_302 (N7229, {N7090_1, N7093});
or_n #(2, 0, 0) OR_138 (N7236, {N7173, N7125});
or_n #(2, 0, 0) OR_139 (N7239, {N7174, N7126});
or_n #(2, 0, 0) OR_140 (N7242, {N7175, N7127});
or_n #(2, 0, 0) OR_141 (N7245, {N7176, N7040});
or_n #(2, 0, 0) OR_142 (N7250, {N7178, N7139});
or_n #(2, 0, 0) OR_143 (N7257, {N7179, N7140});
or_n #(2, 0, 0) OR_144 (N7260, {N7180, N7141});
or_n #(2, 0, 0) OR_145 (N7263, {N7181, N7064});
nand_n #(2, 0, 0) NAND_303 (N7268, {N6792_1, N7183});
nand_n #(2, 0, 0) NAND_304 (N7269, {N6795_1, N7185});
or_n #(3, 0, 0) OR_146 (N7270, {N4957, N7187, N3782});
or_n #(3, 0, 0) OR_147 (N7276, {N4958, N7188, N3783});
or_n #(3, 0, 0) OR_148 (N7282, {N4959, N7189, N3784});
or_n #(3, 0, 0) OR_149 (N7288, {N4961, N7196, N3787});
or_n #(3, 0, 0) OR_150 (N7294, {N3998, N7197, N3788});
nand_n #(2, 0, 0) NAND_305 (N7300, {N7003_1, N7205});
nand_n #(2, 0, 0) NAND_306 (N7301, {N7206, N7151});
or_n #(3, 0, 0) OR_151 (N7304, {N4980, N7207, N3800});
or_n #(3, 0, 0) OR_152 (N7310, {N4984, N7208, N3805});
nand_n #(2, 0, 0) NAND_307 (N7320, {N6891_1, N7215});
nand_n #(2, 0, 0) NAND_308 (N7321, {N6897_1, N7217});
nand_n #(2, 0, 0) NAND_309 (N7328, {N6916_1, N7228});
and_n #(3, 0, 0) AND_583 (N7338, {N7190_0, N1185_6, N2692_1});
and_n #(3, 0, 0) AND_584 (N7339, {N7198_0, N2681_6, N2692_2});
and_n #(3, 0, 0) AND_585 (N7340, {N7190_1, N1247_6, N2767_1});
and_n #(3, 0, 0) AND_586 (N7341, {N7198_1, N2756_6, N2767_2});
and_n #(3, 0, 0) AND_587 (N7342, {N7190_2, N1327_6, N2790_1});
and_n #(3, 0, 0) AND_588 (N7349, {N7198_2, N2779_6, N2790_2});
and_n #(3, 0, 0) AND_589 (N7357, {N7198_3, N2801_6, N2812_1});
notg #(0, 0) NOT_498 (N7363, N7198_4);
and_n #(3, 0, 0) AND_590 (N7364, {N7190_3, N1351_6, N2812_2});
notg #(0, 0) NOT_499 (N7365, N7190_4);
nand_n #(2, 0, 0) NAND_310 (N7394, {N7268, N7184});
nand_n #(2, 0, 0) NAND_311 (N7397, {N7269, N7186});
nand_n #(2, 0, 0) NAND_312 (N7402, {N7204, N7300});
notg #(0, 0) NOT_500 (N7405, N7209_0);
nand_n #(2, 0, 0) NAND_313 (N7406, {N7209_1, N6884});
notg #(0, 0) NOT_501 (N7407, N7212_0);
nand_n #(2, 0, 0) NAND_314 (N7408, {N7212_1, N6888});
nand_n #(2, 0, 0) NAND_315 (N7409, {N7320, N7216});
nand_n #(2, 0, 0) NAND_316 (N7412, {N7321, N7218});
notg #(0, 0) NOT_502 (N7415, N7219_0);
nand_n #(2, 0, 0) NAND_317 (N7416, {N7219_1, N6904});
notg #(0, 0) NOT_503 (N7417, N7222_0);
nand_n #(2, 0, 0) NAND_318 (N7418, {N7222_1, N6908});
notg #(0, 0) NOT_504 (N7419, N7225_0);
nand_n #(2, 0, 0) NAND_319 (N7420, {N7225_1, N6913});
nand_n #(2, 0, 0) NAND_320 (N7421, {N7328, N7229});
notg #(0, 0) NOT_505 (N7424, N7245_0);
notg #(0, 0) NOT_506 (N7425, N7242_0);
notg #(0, 0) NOT_507 (N7426, N7239_0);
notg #(0, 0) NOT_508 (N7427, N7236_0);
notg #(0, 0) NOT_509 (N7428, N7263_0);
notg #(0, 0) NOT_510 (N7429, N7260_0);
notg #(0, 0) NOT_511 (N7430, N7257_0);
notg #(0, 0) NOT_512 (N7431, N7250_0);
notg #(0, 0) NOT_513 (N7432, N7250_1);
and_n #(3, 0, 0) AND_591 (N7433, {N7310_0, N2653_5, N2664_0});
and_n #(3, 0, 0) AND_592 (N7434, {N7304_0, N1161_6, N2664_1});
or_n #(4, 0, 0) OR_153 (N7435, {N7011, N7338, N3621, N2591});
and_n #(3, 0, 0) AND_593 (N7436, {N7270_0, N1185_7, N2692_3});
and_n #(3, 0, 0) AND_594 (N7437, {N7288_0, N2681_7, N2692_4});
and_n #(3, 0, 0) AND_595 (N7438, {N7276_0, N1185_8, N2692_5});
and_n #(3, 0, 0) AND_596 (N7439, {N7294_0, N2681_8, N2692_6});
and_n #(3, 0, 0) AND_597 (N7440, {N7282_0, N1185_9, N2692_7});
and_n #(3, 0, 0) AND_598 (N7441, {N7310_1, N2728_5, N2739_0});
and_n #(3, 0, 0) AND_599 (N7442, {N7304_1, N1223_6, N2739_1});
or_n #(4, 0, 0) OR_154 (N7443, {N7012, N7340, N3632, N2600});
and_n #(3, 0, 0) AND_600 (N7444, {N7270_1, N1247_7, N2767_3});
and_n #(3, 0, 0) AND_601 (N7445, {N7288_1, N2756_7, N2767_4});
and_n #(3, 0, 0) AND_602 (N7446, {N7276_1, N1247_8, N2767_5});
and_n #(3, 0, 0) AND_603 (N7447, {N7294_1, N2756_8, N2767_6});
and_n #(3, 0, 0) AND_604 (N7448, {N7282_1, N1247_9, N2767_7});
or_n #(4, 0, 0) OR_155 (N7449, {N7013, N7342, N3641, N2605});
and_n #(3, 0, 0) AND_605 (N7450, {N7310_2, N3041_5, N3052_0});
and_n #(3, 0, 0) AND_606 (N7451, {N7304_2, N1697_6, N3052_1});
and_n #(3, 0, 0) AND_607 (N7452, {N7294_2, N2779_7, N2790_3});
and_n #(3, 0, 0) AND_608 (N7453, {N7282_2, N1327_7, N2790_4});
and_n #(3, 0, 0) AND_609 (N7454, {N7288_2, N2779_8, N2790_5});
and_n #(3, 0, 0) AND_610 (N7455, {N7276_2, N1327_8, N2790_6});
and_n #(3, 0, 0) AND_611 (N7456, {N7270_2, N1327_9, N2790_7});
and_n #(3, 0, 0) AND_612 (N7457, {N7310_3, N3075_5, N3086_0});
and_n #(3, 0, 0) AND_613 (N7458, {N7304_3, N1731_6, N3086_1});
and_n #(3, 0, 0) AND_614 (N7459, {N7294_3, N2801_7, N2812_3});
and_n #(3, 0, 0) AND_615 (N7460, {N7282_3, N1351_7, N2812_4});
and_n #(3, 0, 0) AND_616 (N7461, {N7288_3, N2801_8, N2812_5});
and_n #(3, 0, 0) AND_617 (N7462, {N7276_3, N1351_8, N2812_6});
and_n #(3, 0, 0) AND_618 (N7463, {N7270_3, N1351_9, N2812_7});
and_n #(3, 0, 0) AND_619 (N7464, {N7250_2, N603_2, N599_2});
notg #(0, 0) NOT_514 (N7465, N7310_4);
notg #(0, 0) NOT_515 (N7466, N7294_4);
notg #(0, 0) NOT_516 (N7467, N7288_4);
notg #(0, 0) NOT_517 (N7468, N7301_0);
or_n #(4, 0, 0) OR_156 (N7469, {N7016, N7364, N3660, N2626});
notg #(0, 0) NOT_518 (N7470, N7304_4);
notg #(0, 0) NOT_519 (N7471, N7282_4);
notg #(0, 0) NOT_520 (N7472, N7276_4);
notg #(0, 0) NOT_521 (N7473, N7270_4);
bufg #(0, 0) BUF_312 (N7474, N7394_0);
bufg #(0, 0) BUF_313 (N7476, N7397_0);
and_n #(2, 0, 0) AND_620 (N7479, {N7301_1, N3068_0});
and_n #(3, 0, 0) AND_621 (N7481, {N7245_1, N1793_2, N3158_6});
and_n #(3, 0, 0) AND_622 (N7482, {N7242_1, N1793_3, N3158_7});
and_n #(3, 0, 0) AND_623 (N7483, {N7239_1, N1793_4, N3158_8});
and_n #(3, 0, 0) AND_624 (N7484, {N7236_1, N1793_5, N3158_9});
and_n #(3, 0, 0) AND_625 (N7485, {N7263_1, N1807_2, N3180_6});
and_n #(3, 0, 0) AND_626 (N7486, {N7260_1, N1807_3, N3180_7});
and_n #(3, 0, 0) AND_627 (N7487, {N7257_1, N1807_4, N3180_8});
and_n #(3, 0, 0) AND_628 (N7488, {N7250_3, N1807_5, N3180_9});
nand_n #(2, 0, 0) NAND_321 (N7489, {N6979_1, N7250_4});
nand_n #(2, 0, 0) NAND_322 (N7492, {N6516_1, N7405});
nand_n #(2, 0, 0) NAND_323 (N7493, {N6526_1, N7407});
nand_n #(2, 0, 0) NAND_324 (N7498, {N6592_1, N7415});
nand_n #(2, 0, 0) NAND_325 (N7499, {N6599_1, N7417});
nand_n #(2, 0, 0) NAND_326 (N7500, {N6609_1, N7419});
and_n #(9, 0, 0) AND_629 (N7503, {N7105, N7166, N7167, N7168, N7169, N7424, N7425, N7426, N7427});
and_n #(9, 0, 0) AND_630 (N7504, {N6640, N7110, N7170, N7171, N7172, N7428, N7429, N7430, N7431});
or_n #(4, 0, 0) OR_157 (N7505, {N7433, N7434, N3616, N2585});
and_n #(2, 0, 0) AND_631 (N7506, {N7435, N2675_0});
or_n #(4, 0, 0) OR_158 (N7507, {N7339, N7436, N3622, N2592});
or_n #(4, 0, 0) OR_159 (N7508, {N7437, N7438, N3623, N2593});
or_n #(4, 0, 0) OR_160 (N7509, {N7439, N7440, N3624, N2594});
or_n #(4, 0, 0) OR_161 (N7510, {N7441, N7442, N3627, N2595});
and_n #(2, 0, 0) AND_632 (N7511, {N7443, N2750_0});
or_n #(4, 0, 0) OR_162 (N7512, {N7341, N7444, N3633, N2601});
or_n #(4, 0, 0) OR_163 (N7513, {N7445, N7446, N3634, N2602});
or_n #(4, 0, 0) OR_164 (N7514, {N7447, N7448, N3635, N2603});
or_n #(4, 0, 0) OR_165 (N7515, {N7450, N7451, N3646, N2610});
or_n #(4, 0, 0) OR_166 (N7516, {N7452, N7453, N3647, N2611});
or_n #(4, 0, 0) OR_167 (N7517, {N7454, N7455, N3648, N2612});
or_n #(4, 0, 0) OR_168 (N7518, {N7349, N7456, N3649, N2613});
or_n #(4, 0, 0) OR_169 (N7519, {N7457, N7458, N3654, N2618});
or_n #(4, 0, 0) OR_170 (N7520, {N7459, N7460, N3655, N2619});
or_n #(4, 0, 0) OR_171 (N7521, {N7461, N7462, N3656, N2620});
or_n #(4, 0, 0) OR_172 (N7522, {N7357, N7463, N3657, N2621});
or_n #(4, 0, 0) OR_173 (N7525, {N4741, N7114, N2624, N7464});
and_n #(3, 0, 0) AND_633 (N7526, {N7468, N3119_9, N3130_8});
notg #(0, 0) NOT_522 (N7527, N7394_1);
notg #(0, 0) NOT_523 (N7528, N7397_1);
notg #(0, 0) NOT_524 (N7529, N7402_0);
and_n #(2, 0, 0) AND_634 (N7530, {N7402_1, N3068_1});
or_n #(3, 0, 0) OR_174 (N7531, {N4981, N7481, N3801});
or_n #(3, 0, 0) OR_175 (N7537, {N4982, N7482, N3802});
or_n #(3, 0, 0) OR_176 (N7543, {N4983, N7483, N3803});
or_n #(3, 0, 0) OR_177 (N7549, {N5165, N7484, N3804});
or_n #(3, 0, 0) OR_178 (N7555, {N4985, N7485, N3806});
or_n #(3, 0, 0) OR_179 (N7561, {N4986, N7486, N3807});
or_n #(3, 0, 0) OR_180 (N7567, {N4547, N7487, N3808});
or_n #(3, 0, 0) OR_181 (N7573, {N4987, N7488, N3809});
nand_n #(2, 0, 0) NAND_327 (N7579, {N7492, N7406});
nand_n #(2, 0, 0) NAND_328 (N7582, {N7493, N7408});
notg #(0, 0) NOT_525 (N7585, N7409_0);
nand_n #(2, 0, 0) NAND_329 (N7586, {N7409_1, N6894});
notg #(0, 0) NOT_526 (N7587, N7412_0);
nand_n #(2, 0, 0) NAND_330 (N7588, {N7412_1, N6900});
nand_n #(2, 0, 0) NAND_331 (N7589, {N7498, N7416});
nand_n #(2, 0, 0) NAND_332 (N7592, {N7499, N7418});
nand_n #(2, 0, 0) NAND_333 (N7595, {N7500, N7420});
notg #(0, 0) NOT_527 (N7598, N7421_0);
nand_n #(2, 0, 0) NAND_334 (N7599, {N7421_1, N6919});
and_n #(2, 0, 0) AND_635 (N7600, {N7505, N2647_0});
and_n #(2, 0, 0) AND_636 (N7601, {N7507, N2675_1});
and_n #(2, 0, 0) AND_637 (N7602, {N7508, N2675_2});
and_n #(2, 0, 0) AND_638 (N7603, {N7509, N2675_3});
and_n #(2, 0, 0) AND_639 (N7604, {N7510, N2722_0});
and_n #(2, 0, 0) AND_640 (N7605, {N7512, N2750_1});
and_n #(2, 0, 0) AND_641 (N7606, {N7513, N2750_2});
and_n #(2, 0, 0) AND_642 (N7607, {N7514, N2750_3});
and_n #(2, 0, 0) AND_643 (N7624, {N6979_2, N7489_0});
and_n #(2, 0, 0) AND_644 (N7625, {N7489_1, N7250_5});
and_n #(2, 0, 0) AND_645 (N7626, {N1149, N7525});
and_n #(5, 0, 0) AND_646 (N7631, {N562_2, N7527, N7528, N6805, N6930});
and_n #(3, 0, 0) AND_647 (N7636, {N7529, N3097_9, N3108_8});
nand_n #(2, 0, 0) NAND_335 (N7657, {N6539_1, N7585});
nand_n #(2, 0, 0) NAND_336 (N7658, {N6556_1, N7587});
nand_n #(2, 0, 0) NAND_337 (N7665, {N6622_1, N7598});
and_n #(3, 0, 0) AND_648 (N7666, {N7555_0, N2653_6, N2664_2});
and_n #(3, 0, 0) AND_649 (N7667, {N7531_0, N1161_7, N2664_3});
and_n #(3, 0, 0) AND_650 (N7668, {N7561_0, N2653_7, N2664_4});
and_n #(3, 0, 0) AND_651 (N7669, {N7537_0, N1161_8, N2664_5});
and_n #(3, 0, 0) AND_652 (N7670, {N7567_0, N2653_8, N2664_6});
and_n #(3, 0, 0) AND_653 (N7671, {N7543_0, N1161_9, N2664_7});
and_n #(3, 0, 0) AND_654 (N7672, {N7573_0, N2653_9, N2664_8});
and_n #(3, 0, 0) AND_655 (N7673, {N7549_0, N1161_10, N2664_9});
and_n #(3, 0, 0) AND_656 (N7674, {N7555_1, N2728_6, N2739_2});
and_n #(3, 0, 0) AND_657 (N7675, {N7531_1, N1223_7, N2739_3});
and_n #(3, 0, 0) AND_658 (N7676, {N7561_1, N2728_7, N2739_4});
and_n #(3, 0, 0) AND_659 (N7677, {N7537_1, N1223_8, N2739_5});
and_n #(3, 0, 0) AND_660 (N7678, {N7567_1, N2728_8, N2739_6});
and_n #(3, 0, 0) AND_661 (N7679, {N7543_1, N1223_9, N2739_7});
and_n #(3, 0, 0) AND_662 (N7680, {N7573_1, N2728_9, N2739_8});
and_n #(3, 0, 0) AND_663 (N7681, {N7549_1, N1223_10, N2739_9});
and_n #(3, 0, 0) AND_664 (N7682, {N7573_2, N3075_6, N3086_2});
and_n #(3, 0, 0) AND_665 (N7683, {N7549_2, N1731_7, N3086_3});
and_n #(3, 0, 0) AND_666 (N7684, {N7573_3, N3041_6, N3052_2});
and_n #(3, 0, 0) AND_667 (N7685, {N7549_3, N1697_7, N3052_3});
and_n #(3, 0, 0) AND_668 (N7686, {N7567_2, N3041_7, N3052_4});
and_n #(3, 0, 0) AND_669 (N7687, {N7543_2, N1697_8, N3052_5});
and_n #(3, 0, 0) AND_670 (N7688, {N7561_2, N3041_8, N3052_6});
and_n #(3, 0, 0) AND_671 (N7689, {N7537_2, N1697_9, N3052_7});
and_n #(3, 0, 0) AND_672 (N7690, {N7555_2, N3041_9, N3052_8});
and_n #(3, 0, 0) AND_673 (N7691, {N7531_2, N1697_10, N3052_9});
and_n #(3, 0, 0) AND_674 (N7692, {N7567_3, N3075_7, N3086_4});
and_n #(3, 0, 0) AND_675 (N7693, {N7543_3, N1731_8, N3086_5});
and_n #(3, 0, 0) AND_676 (N7694, {N7561_3, N3075_8, N3086_6});
and_n #(3, 0, 0) AND_677 (N7695, {N7537_3, N1731_9, N3086_7});
and_n #(3, 0, 0) AND_678 (N7696, {N7555_3, N3075_9, N3086_8});
and_n #(3, 0, 0) AND_679 (N7697, {N7531_3, N1731_10, N3086_9});
or_n #(2, 0, 0) OR_182 (N7698, {N7624, N7625});
notg #(0, 0) NOT_528 (N7699, N7573_4);
notg #(0, 0) NOT_529 (N7700, N7567_4);
notg #(0, 0) NOT_530 (N7701, N7561_4);
notg #(0, 0) NOT_531 (N7702, N7555_4);
and_n #(3, 0, 0) AND_680 (N7703, {N1156, N7631, N245_1});
notg #(0, 0) NOT_532 (N7704, N7549_4);
notg #(0, 0) NOT_533 (N7705, N7543_4);
notg #(0, 0) NOT_534 (N7706, N7537_4);
notg #(0, 0) NOT_535 (N7707, N7531_4);
notg #(0, 0) NOT_536 (N7708, N7579_0);
nand_n #(2, 0, 0) NAND_338 (N7709, {N7579_1, N6739});
notg #(0, 0) NOT_537 (N7710, N7582_0);
nand_n #(2, 0, 0) NAND_339 (N7711, {N7582_1, N6744});
nand_n #(2, 0, 0) NAND_340 (N7712, {N7657, N7586});
nand_n #(2, 0, 0) NAND_341 (N7715, {N7658, N7588});
notg #(0, 0) NOT_538 (N7718, N7589_0);
nand_n #(2, 0, 0) NAND_342 (N7719, {N7589_1, N6772});
notg #(0, 0) NOT_539 (N7720, N7592_0);
nand_n #(2, 0, 0) NAND_343 (N7721, {N7592_1, N6776});
notg #(0, 0) NOT_540 (N7722, N7595_0);
nand_n #(2, 0, 0) NAND_344 (N7723, {N7595_1, N5733});
nand_n #(2, 0, 0) NAND_345 (N7724, {N7665, N7599});
or_n #(4, 0, 0) OR_183 (N7727, {N7666, N7667, N3617, N2586});
or_n #(4, 0, 0) OR_184 (N7728, {N7668, N7669, N3618, N2587});
or_n #(4, 0, 0) OR_185 (N7729, {N7670, N7671, N3619, N2588});
or_n #(4, 0, 0) OR_186 (N7730, {N7672, N7673, N3620, N2589});
or_n #(4, 0, 0) OR_187 (N7731, {N7674, N7675, N3628, N2596});
or_n #(4, 0, 0) OR_188 (N7732, {N7676, N7677, N3629, N2597});
or_n #(4, 0, 0) OR_189 (N7733, {N7678, N7679, N3630, N2598});
or_n #(4, 0, 0) OR_190 (N7734, {N7680, N7681, N3631, N2599});
or_n #(4, 0, 0) OR_191 (N7735, {N7682, N7683, N3638, N2604});
or_n #(4, 0, 0) OR_192 (N7736, {N7684, N7685, N3642, N2606});
or_n #(4, 0, 0) OR_193 (N7737, {N7686, N7687, N3643, N2607});
or_n #(4, 0, 0) OR_194 (N7738, {N7688, N7689, N3644, N2608});
or_n #(4, 0, 0) OR_195 (N7739, {N7690, N7691, N3645, N2609});
or_n #(4, 0, 0) OR_196 (N7740, {N7692, N7693, N3651, N2615});
or_n #(4, 0, 0) OR_197 (N7741, {N7694, N7695, N3652, N2616});
or_n #(4, 0, 0) OR_198 (N7742, {N7696, N7697, N3653, N2617});
nand_n #(2, 0, 0) NAND_346 (N7743, {N6271_1, N7708});
nand_n #(2, 0, 0) NAND_347 (N7744, {N6283_1, N7710});
nand_n #(2, 0, 0) NAND_348 (N7749, {N6341_1, N7718});
nand_n #(2, 0, 0) NAND_349 (N7750, {N6347_1, N7720});
nand_n #(2, 0, 0) NAND_350 (N7751, {N5214_1, N7722});
and_n #(2, 0, 0) AND_681 (N7754, {N7727, N2647_1});
and_n #(2, 0, 0) AND_682 (N7755, {N7728, N2647_2});
and_n #(2, 0, 0) AND_683 (N7756, {N7729, N2647_3});
and_n #(2, 0, 0) AND_684 (N7757, {N7730, N2647_4});
and_n #(2, 0, 0) AND_685 (N7758, {N7731, N2722_1});
and_n #(2, 0, 0) AND_686 (N7759, {N7732, N2722_2});
and_n #(2, 0, 0) AND_687 (N7760, {N7733, N2722_3});
and_n #(2, 0, 0) AND_688 (N7761, {N7734, N2722_4});
nand_n #(2, 0, 0) NAND_351 (N7762, {N7743, N7709});
nand_n #(2, 0, 0) NAND_352 (N7765, {N7744, N7711});
notg #(0, 0) NOT_541 (N7768, N7712_0);
nand_n #(2, 0, 0) NAND_353 (N7769, {N7712_1, N6751});
notg #(0, 0) NOT_542 (N7770, N7715_0);
nand_n #(2, 0, 0) NAND_354 (N7771, {N7715_1, N6760});
nand_n #(2, 0, 0) NAND_355 (N7772, {N7749, N7719});
nand_n #(2, 0, 0) NAND_356 (N7775, {N7750, N7721});
nand_n #(2, 0, 0) NAND_357 (N7778, {N7751, N7723});
notg #(0, 0) NOT_543 (N7781, N7724_0);
nand_n #(2, 0, 0) NAND_358 (N7782, {N7724_1, N5735});
nand_n #(2, 0, 0) NAND_359 (N7787, {N6295_1, N7768});
nand_n #(2, 0, 0) NAND_360 (N7788, {N6313_1, N7770});
nand_n #(2, 0, 0) NAND_361 (N7795, {N5220_1, N7781});
notg #(0, 0) NOT_544 (N7796, N7762_0);
nand_n #(2, 0, 0) NAND_362 (N7797, {N7762_1, N6740});
notg #(0, 0) NOT_545 (N7798, N7765_0);
nand_n #(2, 0, 0) NAND_363 (N7799, {N7765_1, N6745});
nand_n #(2, 0, 0) NAND_364 (N7800, {N7787, N7769});
nand_n #(2, 0, 0) NAND_365 (N7803, {N7788, N7771});
notg #(0, 0) NOT_546 (N7806, N7772_0);
nand_n #(2, 0, 0) NAND_366 (N7807, {N7772_1, N6773});
notg #(0, 0) NOT_547 (N7808, N7775_0);
nand_n #(2, 0, 0) NAND_367 (N7809, {N7775_1, N6777});
notg #(0, 0) NOT_548 (N7810, N7778_0);
nand_n #(2, 0, 0) NAND_368 (N7811, {N7778_1, N6782});
nand_n #(2, 0, 0) NAND_369 (N7812, {N7795, N7782});
nand_n #(2, 0, 0) NAND_370 (N7815, {N6274_1, N7796});
nand_n #(2, 0, 0) NAND_371 (N7816, {N6286_1, N7798});
nand_n #(2, 0, 0) NAND_372 (N7821, {N6344_1, N7806});
nand_n #(2, 0, 0) NAND_373 (N7822, {N6350_1, N7808});
nand_n #(2, 0, 0) NAND_374 (N7823, {N6353_1, N7810});
nand_n #(2, 0, 0) NAND_375 (N7826, {N7815, N7797});
nand_n #(2, 0, 0) NAND_376 (N7829, {N7816, N7799});
notg #(0, 0) NOT_549 (N7832, N7800_0);
nand_n #(2, 0, 0) NAND_377 (N7833, {N7800_1, N6752});
notg #(0, 0) NOT_550 (N7834, N7803_0);
nand_n #(2, 0, 0) NAND_378 (N7835, {N7803_1, N6761});
nand_n #(2, 0, 0) NAND_379 (N7836, {N7821, N7807});
nand_n #(2, 0, 0) NAND_380 (N7839, {N7822, N7809});
nand_n #(2, 0, 0) NAND_381 (N7842, {N7823, N7811});
notg #(0, 0) NOT_551 (N7845, N7812_0);
nand_n #(2, 0, 0) NAND_382 (N7846, {N7812_1, N6790});
nand_n #(2, 0, 0) NAND_383 (N7851, {N6298_1, N7832});
nand_n #(2, 0, 0) NAND_384 (N7852, {N6316_1, N7834});
nand_n #(2, 0, 0) NAND_385 (N7859, {N6364_1, N7845});
notg #(0, 0) NOT_552 (N7860, N7826_0);
nand_n #(2, 0, 0) NAND_386 (N7861, {N7826_1, N6741});
notg #(0, 0) NOT_553 (N7862, N7829_0);
nand_n #(2, 0, 0) NAND_387 (N7863, {N7829_1, N6746});
nand_n #(2, 0, 0) NAND_388 (N7864, {N7851, N7833});
nand_n #(2, 0, 0) NAND_389 (N7867, {N7852, N7835});
notg #(0, 0) NOT_554 (N7870, N7836_0);
nand_n #(2, 0, 0) NAND_390 (N7871, {N7836_1, N5730});
notg #(0, 0) NOT_555 (N7872, N7839_0);
nand_n #(2, 0, 0) NAND_391 (N7873, {N7839_1, N5732});
notg #(0, 0) NOT_556 (N7874, N7842_0);
nand_n #(2, 0, 0) NAND_392 (N7875, {N7842_1, N6783});
nand_n #(2, 0, 0) NAND_393 (N7876, {N7859, N7846});
nand_n #(2, 0, 0) NAND_394 (N7879, {N6277_1, N7860});
nand_n #(2, 0, 0) NAND_395 (N7880, {N6289_1, N7862});
nand_n #(2, 0, 0) NAND_396 (N7885, {N5199_1, N7870});
nand_n #(2, 0, 0) NAND_397 (N7886, {N5208_1, N7872});
nand_n #(2, 0, 0) NAND_398 (N7887, {N6356_1, N7874});
nand_n #(2, 0, 0) NAND_399 (N7890, {N7879, N7861});
nand_n #(2, 0, 0) NAND_400 (N7893, {N7880, N7863});
notg #(0, 0) NOT_557 (N7896, N7864_0);
nand_n #(2, 0, 0) NAND_401 (N7897, {N7864_1, N6753});
notg #(0, 0) NOT_558 (N7898, N7867_0);
nand_n #(2, 0, 0) NAND_402 (N7899, {N7867_1, N6762});
nand_n #(2, 0, 0) NAND_403 (N7900, {N7885, N7871});
nand_n #(2, 0, 0) NAND_404 (N7903, {N7886, N7873});
nand_n #(2, 0, 0) NAND_405 (N7906, {N7887, N7875});
notg #(0, 0) NOT_559 (N7909, N7876_0);
nand_n #(2, 0, 0) NAND_406 (N7910, {N7876_1, N6791});
nand_n #(2, 0, 0) NAND_407 (N7917, {N6301_1, N7896});
nand_n #(2, 0, 0) NAND_408 (N7918, {N6319_1, N7898});
nand_n #(2, 0, 0) NAND_409 (N7923, {N6367_1, N7909});
notg #(0, 0) NOT_560 (N7924, N7890_0);
nand_n #(2, 0, 0) NAND_410 (N7925, {N7890_1, N6680});
notg #(0, 0) NOT_561 (N7926, N7893_0);
nand_n #(2, 0, 0) NAND_411 (N7927, {N7893_1, N6681});
notg #(0, 0) NOT_562 (N7928, N7900_0);
nand_n #(2, 0, 0) NAND_412 (N7929, {N7900_1, N5690});
notg #(0, 0) NOT_563 (N7930, N7903_0);
nand_n #(2, 0, 0) NAND_413 (N7931, {N7903_1, N5691});
nand_n #(2, 0, 0) NAND_414 (N7932, {N7917, N7897});
nand_n #(2, 0, 0) NAND_415 (N7935, {N7918, N7899});
notg #(0, 0) NOT_564 (N7938, N7906_0);
nand_n #(2, 0, 0) NAND_416 (N7939, {N7906_1, N6784});
nand_n #(2, 0, 0) NAND_417 (N7940, {N7923, N7910});
nand_n #(2, 0, 0) NAND_418 (N7943, {N6280_1, N7924});
nand_n #(2, 0, 0) NAND_419 (N7944, {N6292_1, N7926});
nand_n #(2, 0, 0) NAND_420 (N7945, {N5202_1, N7928});
nand_n #(2, 0, 0) NAND_421 (N7946, {N5211_1, N7930});
nand_n #(2, 0, 0) NAND_422 (N7951, {N6359_1, N7938});
nand_n #(2, 0, 0) NAND_423 (N7954, {N7943, N7925});
nand_n #(2, 0, 0) NAND_424 (N7957, {N7944, N7927});
nand_n #(2, 0, 0) NAND_425 (N7960, {N7945, N7929});
nand_n #(2, 0, 0) NAND_426 (N7963, {N7946, N7931});
notg #(0, 0) NOT_565 (N7966, N7932_0);
nand_n #(2, 0, 0) NAND_427 (N7967, {N7932_1, N6754});
notg #(0, 0) NOT_566 (N7968, N7935_0);
nand_n #(2, 0, 0) NAND_428 (N7969, {N7935_1, N6755});
nand_n #(2, 0, 0) NAND_429 (N7970, {N7951, N7939});
notg #(0, 0) NOT_567 (N7973, N7940_0);
nand_n #(2, 0, 0) NAND_430 (N7974, {N7940_1, N6785});
nand_n #(2, 0, 0) NAND_431 (N7984, {N6304_1, N7966});
nand_n #(2, 0, 0) NAND_432 (N7985, {N6322_1, N7968});
nand_n #(2, 0, 0) NAND_433 (N7987, {N6370_1, N7973});
and_n #(3, 0, 0) AND_689 (N7988, {N7957_0, N6831_1, N1157_0});
and_n #(3, 0, 0) AND_690 (N7989, {N7954_0, N6415_2, N1157_1});
and_n #(3, 0, 0) AND_691 (N7990, {N7957_1, N7041_1, N566_1});
and_n #(3, 0, 0) AND_692 (N7991, {N7954_1, N7177, N566_2});
notg #(0, 0) NOT_568 (N7992, N7970_0);
nand_n #(2, 0, 0) NAND_434 (N7993, {N7970_1, N6448});
and_n #(3, 0, 0) AND_693 (N7994, {N7963_0, N6857_1, N1219_0});
and_n #(3, 0, 0) AND_694 (N7995, {N7960_0, N6441_2, N1219_1});
and_n #(3, 0, 0) AND_695 (N7996, {N7963_1, N7065_1, N583_1});
and_n #(3, 0, 0) AND_696 (N7997, {N7960_1, N7182, N583_2});
nand_n #(2, 0, 0) NAND_435 (N7998, {N7984, N7967});
nand_n #(2, 0, 0) NAND_436 (N8001, {N7985, N7969});
nand_n #(2, 0, 0) NAND_437 (N8004, {N7987, N7974});
nand_n #(2, 0, 0) NAND_438 (N8009, {N6051_1, N7992});
or_n #(4, 0, 0) OR_199 (N8013, {N7988, N7989, N7990, N7991});
or_n #(4, 0, 0) OR_200 (N8017, {N7994, N7995, N7996, N7997});
notg #(0, 0) NOT_569 (N8020, N7998_0);
nand_n #(2, 0, 0) NAND_439 (N8021, {N7998_1, N6682});
notg #(0, 0) NOT_570 (N8022, N8001_0);
nand_n #(2, 0, 0) NAND_440 (N8023, {N8001_1, N6683});
nand_n #(2, 0, 0) NAND_441 (N8025, {N8009, N7993});
notg #(0, 0) NOT_571 (N8026, N8004_0);
nand_n #(2, 0, 0) NAND_442 (N8027, {N8004_1, N6449});
nand_n #(2, 0, 0) NAND_443 (N8031, {N6307_1, N8020});
nand_n #(2, 0, 0) NAND_444 (N8032, {N6310_1, N8022});
notg #(0, 0) NOT_572 (N8033, N8013_0);
nand_n #(2, 0, 0) NAND_445 (N8034, {N6054_1, N8026});
and_n #(2, 0, 0) AND_697 (N8035, {N583_3, N8025});
notg #(0, 0) NOT_573 (N8036, N8017_0);
nand_n #(2, 0, 0) NAND_446 (N8037, {N8031, N8021});
nand_n #(2, 0, 0) NAND_447 (N8038, {N8032, N8023});
nand_n #(2, 0, 0) NAND_448 (N8039, {N8034, N8027});
notg #(0, 0) NOT_574 (N8040, N8038);
and_n #(2, 0, 0) AND_698 (N8041, {N566_3, N8037});
notg #(0, 0) NOT_575 (N8042, N8039);
and_n #(2, 0, 0) AND_699 (N8043, {N8040, N1157_2});
and_n #(2, 0, 0) AND_700 (N8044, {N8042, N1219_2});
or_n #(2, 0, 0) OR_201 (N8045, {N8043, N8041});
or_n #(2, 0, 0) OR_202 (N8048, {N8044, N8035});
nand_n #(2, 0, 0) NAND_449 (N8055, {N8045_0, N8033});
notg #(0, 0) NOT_576 (N8056, N8045_1);
nand_n #(2, 0, 0) NAND_450 (N8057, {N8048_0, N8036});
notg #(0, 0) NOT_577 (N8058, N8048_1);
nand_n #(2, 0, 0) NAND_451 (N8059, {N8013_1, N8056});
nand_n #(2, 0, 0) NAND_452 (N8060, {N8017_1, N8058});
nand_n #(2, 0, 0) NAND_453 (N8061, {N8055, N8059});
nand_n #(2, 0, 0) NAND_454 (N8064, {N8057, N8060});
and_n #(3, 0, 0) AND_701 (N8071, {N8064_0, N1777_6, N3130_9});
and_n #(3, 0, 0) AND_702 (N8072, {N8061_0, N1761_6, N3108_9});
notg #(0, 0) NOT_578 (N8073, N8061_1);
notg #(0, 0) NOT_579 (N8074, N8064_1);
or_n #(4, 0, 0) OR_203 (N8075, {N7526, N8071, N3659, N2625});
or_n #(4, 0, 0) OR_204 (N8076, {N7636, N8072, N3661, N2627});
and_n #(2, 0, 0) AND_703 (N8077, {N8073, N1727_1});
and_n #(2, 0, 0) AND_704 (N8078, {N8074, N1727_2});
or_n #(2, 0, 0) OR_205 (N8079, {N7530, N8077});
or_n #(2, 0, 0) OR_206 (N8082, {N7479, N8078});
and_n #(2, 0, 0) AND_705 (N8089, {N8079_0, N3063_0});
and_n #(2, 0, 0) AND_706 (N8090, {N8082_0, N3063_1});
and_n #(2, 0, 0) AND_707 (N8091, {N8079_1, N3063_2});
and_n #(2, 0, 0) AND_708 (N8092, {N8082_1, N3063_3});
or_n #(2, 0, 0) OR_207 (N8093, {N8089, N3071});
or_n #(2, 0, 0) OR_208 (N8096, {N8090, N3072});
or_n #(2, 0, 0) OR_209 (N8099, {N8091, N3073});
or_n #(2, 0, 0) OR_210 (N8102, {N8092, N3074});
and_n #(3, 0, 0) AND_709 (N8113, {N8102_0, N2779_9, N2790_8});
and_n #(3, 0, 0) AND_710 (N8114, {N8099_0, N1327_10, N2790_9});
and_n #(3, 0, 0) AND_711 (N8115, {N8102_1, N2801_9, N2812_8});
and_n #(3, 0, 0) AND_712 (N8116, {N8099_1, N1351_10, N2812_9});
and_n #(3, 0, 0) AND_713 (N8117, {N8096_0, N2681_9, N2692_8});
and_n #(3, 0, 0) AND_714 (N8118, {N8093_0, N1185_10, N2692_9});
and_n #(3, 0, 0) AND_715 (N8119, {N8096_1, N2756_9, N2767_8});
and_n #(3, 0, 0) AND_716 (N8120, {N8093_1, N1247_10, N2767_9});
or_n #(4, 0, 0) OR_211 (N8121, {N8117, N8118, N3662, N2703});
or_n #(4, 0, 0) OR_212 (N8122, {N8119, N8120, N3663, N2778});
or_n #(4, 0, 0) OR_213 (N8123, {N8113, N8114, N3650, N2614});
or_n #(4, 0, 0) OR_214 (N8124, {N8115, N8116, N3658, N2622});
and_n #(2, 0, 0) AND_717 (N8125, {N8121, N2675_4});
and_n #(2, 0, 0) AND_718 (N8126, {N8122, N2750_4});
notg #(0, 0) NOT_580 (N8127, N8125);
notg #(0, 0) NOT_581 (N8128, N8126);

endmodule
