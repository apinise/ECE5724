module c5315 (N1,N4,N11,N14,N17,N20,N23,N24,N25,N26,
              N27,N31,N34,N37,N40,N43,N46,N49,N52,N53,
              N54,N61,N64,N67,N70,N73,N76,N79,N80,N81,
              N82,N83,N86,N87,N88,N91,N94,N97,N100,N103,
              N106,N109,N112,N113,N114,N115,N116,N117,N118,N119,
              N120,N121,N122,N123,N126,N127,N128,N129,N130,N131,
              N132,N135,N136,N137,N140,N141,N145,N146,N149,N152,
              N155,N158,N161,N164,N167,N170,N173,N176,N179,N182,
              N185,N188,N191,N194,N197,N200,N203,N206,N209,N210,
              N217,N218,N225,N226,N233,N234,N241,N242,N245,N248,
              N251,N254,N257,N264,N265,N272,N273,N280,N281,N288,
              N289,N292,N293,N299,N302,N307,N308,N315,N316,N323,
              N324,N331,N332,N335,N338,N341,N348,N351,N358,N361,
              N366,N369,N372,N373,N374,N386,N389,N400,N411,N422,
              N435,N446,N457,N468,N479,N490,N503,N514,N523,N534,
              N545,N549,N552,N556,N559,N562,N566,N571,N574,N577,
              N580,N583,N588,N591,N592,N595,N596,N597,N598,N599,
              N603,N607,N610,N613,N616,N619,N625,N631,N709,N816,
              N1066,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,N1145,
              N1147,N1152,N1153,N1154,N1155,N1972,N2054,N2060,N2061,N2139,
              N2142,N2309,N2387,N2527,N2584,N2590,N2623,N3357,N3358,N3359,
              N3360,N3604,N3613,N4272,N4275,N4278,N4279,N4737,N4738,N4739,
              N4740,N5240,N5388,N6641,N6643,N6646,N6648,N6716,N6877,N6924,
              N6925,N6926,N6927,N7015,N7363,N7365,N7432,N7449,N7465,N7466,
              N7467,N7469,N7470,N7471,N7472,N7473,N7474,N7476,N7503,N7504,
              N7506,N7511,N7515,N7516,N7517,N7518,N7519,N7520,N7521,N7522,
              N7600,N7601,N7602,N7603,N7604,N7605,N7606,N7607,N7626,N7698,
              N7699,N7700,N7701,N7702,N7703,N7704,N7705,N7706,N7707,N7735,
              N7736,N7737,N7738,N7739,N7740,N7741,N7742,N7754,N7755,N7756,
              N7757,N7758,N7759,N7760,N7761,N8075,N8076,N8123,N8124,N8127,
              N8128);

input N1,N4,N11,N14,N17,N20,N23,N24,N25,N26,
      N27,N31,N34,N37,N40,N43,N46,N49,N52,N53,
      N54,N61,N64,N67,N70,N73,N76,N79,N80,N81,
      N82,N83,N86,N87,N88,N91,N94,N97,N100,N103,
      N106,N109,N112,N113,N114,N115,N116,N117,N118,N119,
      N120,N121,N122,N123,N126,N127,N128,N129,N130,N131,
      N132,N135,N136,N137,N140,N141,N145,N146,N149,N152,
      N155,N158,N161,N164,N167,N170,N173,N176,N179,N182,
      N185,N188,N191,N194,N197,N200,N203,N206,N209,N210,
      N217,N218,N225,N226,N233,N234,N241,N242,N245,N248,
      N251,N254,N257,N264,N265,N272,N273,N280,N281,N288,
      N289,N292,N293,N299,N302,N307,N308,N315,N316,N323,
      N324,N331,N332,N335,N338,N341,N348,N351,N358,N361,
      N366,N369,N372,N373,N374,N386,N389,N400,N411,N422,
      N435,N446,N457,N468,N479,N490,N503,N514,N523,N534,
      N545,N549,N552,N556,N559,N562,N566,N571,N574,N577,
      N580,N583,N588,N591,N592,N595,N596,N597,N598,N599,
      N603,N607,N610,N613,N616,N619,N625,N631;

output N709,N816,N1066,N1137,N1138,N1139,N1140,N1141,N1142,N1143,
       N1144,N1145,N1147,N1152,N1153,N1154,N1155,N1972,N2054,N2060,
       N2061,N2139,N2142,N2309,N2387,N2527,N2584,N2590,N2623,N3357,
       N3358,N3359,N3360,N3604,N3613,N4272,N4275,N4278,N4279,N4737,
       N4738,N4739,N4740,N5240,N5388,N6641,N6643,N6646,N6648,N6716,
       N6877,N6924,N6925,N6926,N6927,N7015,N7363,N7365,N7432,N7449,
       N7465,N7466,N7467,N7469,N7470,N7471,N7472,N7473,N7474,N7476,
       N7503,N7504,N7506,N7511,N7515,N7516,N7517,N7518,N7519,N7520,
       N7521,N7522,N7600,N7601,N7602,N7603,N7604,N7605,N7606,N7607,
       N7626,N7698,N7699,N7700,N7701,N7702,N7703,N7704,N7705,N7706,
       N7707,N7735,N7736,N7737,N7738,N7739,N7740,N7741,N7742,N7754,
       N7755,N7756,N7757,N7758,N7759,N7760,N7761,N8075,N8076,N8123,
       N8124,N8127,N8128;

wire N1042,N1043,N1067,N1080,N1092,N1104,N1146,N1148,N1149,N1150,
     N1151,N1156,N1157,N1161,N1173,N1185,N1197,N1209,N1213,N1216,
     N1219,N1223,N1235,N1247,N1259,N1271,N1280,N1292,N1303,N1315,
     N1327,N1339,N1351,N1363,N1375,N1378,N1381,N1384,N1387,N1390,
     N1393,N1396,N1415,N1418,N1421,N1424,N1427,N1430,N1433,N1436,
     N1455,N1462,N1469,N1475,N1479,N1482,N1492,N1495,N1498,N1501,
     N1504,N1507,N1510,N1513,N1516,N1519,N1522,N1525,N1542,N1545,
     N1548,N1551,N1554,N1557,N1560,N1563,N1566,N1573,N1580,N1583,
     N1588,N1594,N1597,N1600,N1603,N1606,N1609,N1612,N1615,N1618,
     N1621,N1624,N1627,N1630,N1633,N1636,N1639,N1642,N1645,N1648,
     N1651,N1654,N1657,N1660,N1663,N1675,N1685,N1697,N1709,N1721,
     N1727,N1731,N1743,N1755,N1758,N1761,N1769,N1777,N1785,N1793,
     N1800,N1807,N1814,N1821,N1824,N1827,N1830,N1833,N1836,N1839,
     N1842,N1845,N1848,N1851,N1854,N1857,N1860,N1863,N1866,N1869,
     N1872,N1875,N1878,N1881,N1884,N1887,N1890,N1893,N1896,N1899,
     N1902,N1905,N1908,N1911,N1914,N1917,N1920,N1923,N1926,N1929,
     N1932,N1935,N1938,N1941,N1944,N1947,N1950,N1953,N1956,N1959,
     N1962,N1965,N1968,N2349,N2350,N2585,N2586,N2587,N2588,N2589,
     N2591,N2592,N2593,N2594,N2595,N2596,N2597,N2598,N2599,N2600,
     N2601,N2602,N2603,N2604,N2605,N2606,N2607,N2608,N2609,N2610,
     N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,N2620,
     N2621,N2622,N2624,N2625,N2626,N2627,N2628,N2629,N2630,N2631,
     N2632,N2633,N2634,N2635,N2636,N2637,N2638,N2639,N2640,N2641,
     N2642,N2643,N2644,N2645,N2646,N2647,N2653,N2664,N2675,N2681,
     N2692,N2703,N2704,N2709,N2710,N2711,N2712,N2713,N2714,N2715,
     N2716,N2717,N2718,N2719,N2720,N2721,N2722,N2728,N2739,N2750,
     N2756,N2767,N2778,N2779,N2790,N2801,N2812,N2823,N2824,N2825,
     N2826,N2827,N2828,N2829,N2830,N2831,N2832,N2833,N2834,N2835,
     N2836,N2837,N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,
     N2846,N2847,N2848,N2849,N2850,N2851,N2852,N2853,N2854,N2855,
     N2861,N2867,N2868,N2869,N2870,N2871,N2872,N2873,N2874,N2875,
     N2876,N2877,N2882,N2891,N2901,N2902,N2903,N2904,N2905,N2906,
     N2907,N2908,N2909,N2910,N2911,N2912,N2913,N2914,N2915,N2916,
     N2917,N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,
     N2927,N2928,N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,
     N2937,N2938,N2939,N2940,N2941,N2942,N2948,N2954,N2955,N2956,
     N2957,N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2969,N2970,
     N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,N2979,N2980,
     N2981,N2982,N2983,N2984,N2985,N2986,N2987,N2988,N2989,N2990,
     N2991,N2992,N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,
     N3003,N3006,N3007,N3010,N3013,N3014,N3015,N3016,N3017,N3018,
     N3019,N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,
     N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3038,N3041,N3052,
     N3063,N3068,N3071,N3072,N3073,N3074,N3075,N3086,N3097,N3108,
     N3119,N3130,N3141,N3142,N3143,N3144,N3145,N3146,N3147,N3158,
     N3169,N3180,N3191,N3194,N3195,N3196,N3197,N3198,N3199,N3200,
     N3203,N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3408,N3409,
     N3410,N3411,N3412,N3413,N3414,N3415,N3416,N3444,N3445,N3446,
     N3447,N3448,N3449,N3450,N3451,N3452,N3453,N3454,N3455,N3456,
     N3459,N3460,N3461,N3462,N3463,N3464,N3465,N3466,N3481,N3482,
     N3483,N3484,N3485,N3486,N3487,N3488,N3489,N3490,N3491,N3492,
     N3493,N3502,N3503,N3504,N3505,N3506,N3507,N3508,N3509,N3510,
     N3511,N3512,N3513,N3514,N3515,N3558,N3559,N3560,N3561,N3562,
     N3563,N3605,N3606,N3607,N3608,N3609,N3610,N3614,N3615,N3616,
     N3617,N3618,N3619,N3620,N3621,N3622,N3623,N3624,N3625,N3626,
     N3627,N3628,N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3636,
     N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,N3646,
     N3647,N3648,N3649,N3650,N3651,N3652,N3653,N3654,N3655,N3656,
     N3657,N3658,N3659,N3660,N3661,N3662,N3663,N3664,N3665,N3666,
     N3667,N3668,N3669,N3670,N3671,N3672,N3673,N3674,N3675,N3676,
     N3677,N3678,N3679,N3680,N3681,N3682,N3683,N3684,N3685,N3686,
     N3687,N3688,N3689,N3691,N3700,N3701,N3702,N3703,N3704,N3705,
     N3708,N3709,N3710,N3711,N3712,N3713,N3715,N3716,N3717,N3718,
     N3719,N3720,N3721,N3722,N3723,N3724,N3725,N3726,N3727,N3728,
     N3729,N3730,N3731,N3732,N3738,N3739,N3740,N3741,N3742,N3743,
     N3744,N3745,N3746,N3747,N3748,N3749,N3750,N3751,N3752,N3753,
     N3754,N3755,N3756,N3757,N3758,N3759,N3760,N3761,N3762,N3763,
     N3764,N3765,N3766,N3767,N3768,N3769,N3770,N3771,N3775,N3779,
     N3780,N3781,N3782,N3783,N3784,N3785,N3786,N3787,N3788,N3789,
     N3793,N3797,N3800,N3801,N3802,N3803,N3804,N3805,N3806,N3807,
     N3808,N3809,N3810,N3813,N3816,N3819,N3822,N3823,N3824,N3827,
     N3828,N3829,N3830,N3831,N3834,N3835,N3836,N3837,N3838,N3839,
     N3840,N3841,N3842,N3849,N3855,N3861,N3867,N3873,N3881,N3887,
     N3893,N3908,N3909,N3911,N3914,N3915,N3916,N3917,N3918,N3919,
     N3920,N3921,N3927,N3933,N3942,N3948,N3956,N3962,N3968,N3975,
     N3976,N3977,N3978,N3979,N3980,N3981,N3982,N3983,N3984,N3987,
     N3988,N3989,N3990,N3991,N3998,N4008,N4011,N4021,N4024,N4027,
     N4031,N4032,N4033,N4034,N4035,N4036,N4037,N4038,N4039,N4040,
     N4041,N4042,N4067,N4080,N4088,N4091,N4094,N4097,N4100,N4103,
     N4106,N4109,N4144,N4147,N4150,N4153,N4156,N4159,N4183,N4184,
     N4185,N4186,N4188,N4191,N4196,N4197,N4198,N4199,N4200,N4203,
     N4206,N4209,N4212,N4215,N4219,N4223,N4224,N4225,N4228,N4231,
     N4234,N4237,N4240,N4243,N4246,N4249,N4252,N4255,N4258,N4263,
     N4264,N4267,N4268,N4269,N4270,N4271,N4273,N4274,N4276,N4277,
     N4280,N4284,N4290,N4297,N4298,N4301,N4305,N4310,N4316,N4320,
     N4325,N4331,N4332,N4336,N4342,N4349,N4357,N4364,N4375,N4379,
     N4385,N4392,N4396,N4400,N4405,N4412,N4418,N4425,N4436,N4440,
     N4445,N4451,N4456,N4462,N4469,N4477,N4512,N4515,N4516,N4521,
     N4523,N4524,N4532,N4547,N4548,N4551,N4554,N4557,N4560,N4563,
     N4566,N4569,N4572,N4575,N4578,N4581,N4584,N4587,N4590,N4593,
     N4596,N4599,N4602,N4605,N4608,N4611,N4614,N4617,N4621,N4624,
     N4627,N4630,N4633,N4637,N4640,N4643,N4646,N4649,N4652,N4655,
     N4658,N4662,N4665,N4668,N4671,N4674,N4677,N4680,N4683,N4686,
     N4689,N4692,N4695,N4698,N4701,N4702,N4720,N4721,N4724,N4725,
     N4726,N4727,N4728,N4729,N4730,N4731,N4732,N4733,N4734,N4735,
     N4736,N4741,N4855,N4856,N4908,N4909,N4939,N4942,N4947,N4953,
     N4954,N4955,N4956,N4957,N4958,N4959,N4960,N4961,N4965,N4966,
     N4967,N4968,N4972,N4973,N4974,N4975,N4976,N4977,N4978,N4979,
     N4980,N4981,N4982,N4983,N4984,N4985,N4986,N4987,N5049,N5052,
     N5053,N5054,N5055,N5056,N5057,N5058,N5059,N5060,N5061,N5062,
     N5063,N5065,N5066,N5067,N5068,N5069,N5070,N5071,N5072,N5073,
     N5074,N5075,N5076,N5077,N5078,N5079,N5080,N5081,N5082,N5083,
     N5084,N5085,N5086,N5087,N5088,N5089,N5090,N5091,N5092,N5093,
     N5094,N5095,N5096,N5097,N5098,N5099,N5100,N5101,N5102,N5103,
     N5104,N5105,N5106,N5107,N5108,N5109,N5110,N5111,N5112,N5113,
     N5114,N5115,N5116,N5117,N5118,N5119,N5120,N5121,N5122,N5123,
     N5124,N5125,N5126,N5127,N5128,N5129,N5130,N5131,N5132,N5133,
     N5135,N5136,N5137,N5138,N5139,N5140,N5141,N5142,N5143,N5144,
     N5145,N5146,N5147,N5148,N5150,N5153,N5154,N5155,N5156,N5157,
     N5160,N5161,N5162,N5163,N5164,N5165,N5166,N5169,N5172,N5173,
     N5176,N5177,N5180,N5183,N5186,N5189,N5192,N5195,N5198,N5199,
     N5202,N5205,N5208,N5211,N5214,N5217,N5220,N5223,N5224,N5225,
     N5226,N5227,N5228,N5229,N5230,N5232,N5233,N5234,N5235,N5236,
     N5239,N5241,N5242,N5243,N5244,N5245,N5246,N5247,N5248,N5249,
     N5250,N5252,N5253,N5254,N5255,N5256,N5257,N5258,N5259,N5260,
     N5261,N5262,N5263,N5264,N5274,N5275,N5282,N5283,N5284,N5298,
     N5299,N5300,N5303,N5304,N5305,N5306,N5307,N5308,N5309,N5310,
     N5311,N5312,N5315,N5319,N5324,N5328,N5331,N5332,N5346,N5363,
     N5364,N5365,N5366,N5367,N5368,N5369,N5370,N5371,N5374,N5377,
     N5382,N5385,N5389,N5396,N5407,N5418,N5424,N5431,N5441,N5452,
     N5462,N5469,N5470,N5477,N5488,N5498,N5506,N5520,N5536,N5549,
     N5555,N5562,N5573,N5579,N5595,N5606,N5616,N5617,N5618,N5619,
     N5620,N5621,N5622,N5624,N5634,N5655,N5671,N5684,N5690,N5691,
     N5692,N5696,N5700,N5703,N5707,N5711,N5726,N5727,N5728,N5730,
     N5731,N5732,N5733,N5734,N5735,N5736,N5739,N5742,N5745,N5755,
     N5756,N5954,N5955,N5956,N6005,N6006,N6023,N6024,N6025,N6028,
     N6031,N6034,N6037,N6040,N6044,N6045,N6048,N6051,N6054,N6065,
     N6066,N6067,N6068,N6069,N6071,N6072,N6073,N6074,N6075,N6076,
     N6077,N6078,N6079,N6080,N6083,N6084,N6085,N6086,N6087,N6088,
     N6089,N6090,N6091,N6094,N6095,N6096,N6097,N6098,N6099,N6100,
     N6101,N6102,N6103,N6104,N6105,N6106,N6107,N6108,N6111,N6112,
     N6113,N6114,N6115,N6116,N6117,N6120,N6121,N6122,N6123,N6124,
     N6125,N6126,N6127,N6128,N6129,N6130,N6131,N6132,N6133,N6134,
     N6135,N6136,N6137,N6138,N6139,N6140,N6143,N6144,N6145,N6146,
     N6147,N6148,N6149,N6152,N6153,N6154,N6155,N6156,N6157,N6158,
     N6159,N6160,N6161,N6162,N6163,N6164,N6168,N6171,N6172,N6173,
     N6174,N6175,N6178,N6179,N6180,N6181,N6182,N6183,N6184,N6185,
     N6186,N6187,N6188,N6189,N6190,N6191,N6192,N6193,N6194,N6197,
     N6200,N6203,N6206,N6209,N6212,N6215,N6218,N6221,N6234,N6235,
     N6238,N6241,N6244,N6247,N6250,N6253,N6256,N6259,N6262,N6265,
     N6268,N6271,N6274,N6277,N6280,N6283,N6286,N6289,N6292,N6295,
     N6298,N6301,N6304,N6307,N6310,N6313,N6316,N6319,N6322,N6325,
     N6328,N6331,N6335,N6338,N6341,N6344,N6347,N6350,N6353,N6356,
     N6359,N6364,N6367,N6370,N6373,N6374,N6375,N6376,N6377,N6378,
     N6382,N6386,N6388,N6392,N6397,N6411,N6415,N6419,N6427,N6434,
     N6437,N6441,N6445,N6448,N6449,N6466,N6469,N6470,N6471,N6472,
     N6473,N6474,N6475,N6476,N6477,N6478,N6482,N6486,N6490,N6494,
     N6500,N6504,N6508,N6512,N6516,N6526,N6536,N6539,N6553,N6556,
     N6566,N6569,N6572,N6575,N6580,N6584,N6587,N6592,N6599,N6606,
     N6609,N6619,N6622,N6630,N6631,N6632,N6633,N6634,N6637,N6640,
     N6650,N6651,N6653,N6655,N6657,N6659,N6660,N6661,N6662,N6663,
     N6664,N6666,N6668,N6670,N6672,N6675,N6680,N6681,N6682,N6683,
     N6689,N6690,N6691,N6692,N6693,N6695,N6698,N6699,N6700,N6703,
     N6708,N6709,N6710,N6711,N6712,N6713,N6714,N6715,N6718,N6719,
     N6720,N6721,N6722,N6724,N6739,N6740,N6741,N6744,N6745,N6746,
     N6751,N6752,N6753,N6754,N6755,N6760,N6761,N6762,N6772,N6773,
     N6776,N6777,N6782,N6783,N6784,N6785,N6790,N6791,N6792,N6795,
     N6801,N6802,N6803,N6804,N6805,N6806,N6807,N6808,N6809,N6810,
     N6811,N6812,N6813,N6814,N6815,N6816,N6817,N6823,N6824,N6825,
     N6826,N6827,N6828,N6829,N6830,N6831,N6834,N6835,N6836,N6837,
     N6838,N6839,N6840,N6841,N6842,N6843,N6844,N6850,N6851,N6852,
     N6853,N6854,N6855,N6856,N6857,N6860,N6861,N6862,N6863,N6866,
     N6872,N6873,N6874,N6875,N6876,N6879,N6880,N6881,N6884,N6885,
     N6888,N6889,N6890,N6891,N6894,N6895,N6896,N6897,N6900,N6901,
     N6904,N6905,N6908,N6909,N6912,N6913,N6914,N6915,N6916,N6919,
     N6922,N6923,N6930,N6932,N6935,N6936,N6937,N6938,N6939,N6940,
     N6946,N6947,N6948,N6949,N6953,N6954,N6955,N6956,N6957,N6958,
     N6964,N6965,N6966,N6967,N6973,N6974,N6975,N6976,N6977,N6978,
     N6979,N6987,N6990,N6999,N7002,N7003,N7006,N7011,N7012,N7013,
     N7016,N7018,N7019,N7020,N7021,N7022,N7023,N7028,N7031,N7034,
     N7037,N7040,N7041,N7044,N7045,N7046,N7047,N7048,N7049,N7054,
     N7057,N7060,N7064,N7065,N7072,N7073,N7074,N7075,N7076,N7079,
     N7080,N7083,N7084,N7085,N7086,N7087,N7088,N7089,N7090,N7093,
     N7094,N7097,N7101,N7105,N7110,N7114,N7115,N7116,N7125,N7126,
     N7127,N7130,N7131,N7139,N7140,N7141,N7146,N7147,N7149,N7150,
     N7151,N7152,N7153,N7158,N7159,N7160,N7166,N7167,N7168,N7169,
     N7170,N7171,N7172,N7173,N7174,N7175,N7176,N7177,N7178,N7179,
     N7180,N7181,N7182,N7183,N7184,N7185,N7186,N7187,N7188,N7189,
     N7190,N7196,N7197,N7198,N7204,N7205,N7206,N7207,N7208,N7209,
     N7212,N7215,N7216,N7217,N7218,N7219,N7222,N7225,N7228,N7229,
     N7236,N7239,N7242,N7245,N7250,N7257,N7260,N7263,N7268,N7269,
     N7270,N7276,N7282,N7288,N7294,N7300,N7301,N7304,N7310,N7320,
     N7321,N7328,N7338,N7339,N7340,N7341,N7342,N7349,N7357,N7364,
     N7394,N7397,N7402,N7405,N7406,N7407,N7408,N7409,N7412,N7415,
     N7416,N7417,N7418,N7419,N7420,N7421,N7424,N7425,N7426,N7427,
     N7428,N7429,N7430,N7431,N7433,N7434,N7435,N7436,N7437,N7438,
     N7439,N7440,N7441,N7442,N7443,N7444,N7445,N7446,N7447,N7448,
     N7450,N7451,N7452,N7453,N7454,N7455,N7456,N7457,N7458,N7459,
     N7460,N7461,N7462,N7463,N7464,N7468,N7479,N7481,N7482,N7483,
     N7484,N7485,N7486,N7487,N7488,N7489,N7492,N7493,N7498,N7499,
     N7500,N7505,N7507,N7508,N7509,N7510,N7512,N7513,N7514,N7525,
     N7526,N7527,N7528,N7529,N7530,N7531,N7537,N7543,N7549,N7555,
     N7561,N7567,N7573,N7579,N7582,N7585,N7586,N7587,N7588,N7589,
     N7592,N7595,N7598,N7599,N7624,N7625,N7631,N7636,N7657,N7658,
     N7665,N7666,N7667,N7668,N7669,N7670,N7671,N7672,N7673,N7674,
     N7675,N7676,N7677,N7678,N7679,N7680,N7681,N7682,N7683,N7684,
     N7685,N7686,N7687,N7688,N7689,N7690,N7691,N7692,N7693,N7694,
     N7695,N7696,N7697,N7708,N7709,N7710,N7711,N7712,N7715,N7718,
     N7719,N7720,N7721,N7722,N7723,N7724,N7727,N7728,N7729,N7730,
     N7731,N7732,N7733,N7734,N7743,N7744,N7749,N7750,N7751,N7762,
     N7765,N7768,N7769,N7770,N7771,N7772,N7775,N7778,N7781,N7782,
     N7787,N7788,N7795,N7796,N7797,N7798,N7799,N7800,N7803,N7806,
     N7807,N7808,N7809,N7810,N7811,N7812,N7815,N7816,N7821,N7822,
     N7823,N7826,N7829,N7832,N7833,N7834,N7835,N7836,N7839,N7842,
     N7845,N7846,N7851,N7852,N7859,N7860,N7861,N7862,N7863,N7864,
     N7867,N7870,N7871,N7872,N7873,N7874,N7875,N7876,N7879,N7880,
     N7885,N7886,N7887,N7890,N7893,N7896,N7897,N7898,N7899,N7900,
     N7903,N7906,N7909,N7910,N7917,N7918,N7923,N7924,N7925,N7926,
     N7927,N7928,N7929,N7930,N7931,N7932,N7935,N7938,N7939,N7940,
     N7943,N7944,N7945,N7946,N7951,N7954,N7957,N7960,N7963,N7966,
     N7967,N7968,N7969,N7970,N7973,N7974,N7984,N7985,N7987,N7988,
     N7989,N7990,N7991,N7992,N7993,N7994,N7995,N7996,N7997,N7998,
     N8001,N8004,N8009,N8013,N8017,N8020,N8021,N8022,N8023,N8025,
     N8026,N8027,N8031,N8032,N8033,N8034,N8035,N8036,N8037,N8038,
     N8039,N8040,N8041,N8042,N8043,N8044,N8045,N8048,N8055,N8056,
     N8057,N8058,N8059,N8060,N8061,N8064,N8071,N8072,N8073,N8074,
     N8077,N8078,N8079,N8082,N8089,N8090,N8091,N8092,N8093,N8096,
     N8099,N8102,N8113,N8114,N8115,N8116,N8117,N8118,N8119,N8120,
     N8121,N8122,N8125,N8126;

buf_1 U178 ( .Z(N709), .A(N141) );
buf_1 U179 ( .Z(N816), .A(N293) );
and2_1 U180 ( .Z(N1042), .A(N135), .B(N631) );
inv_1 U181 ( .Z(N1043), .A(N591) );
buf_1 U182 ( .Z(N1066), .A(N592) );
inv_1 U183 ( .Z(N1067), .A(N595) );
inv_1 U184 ( .Z(N1080), .A(N596) );
inv_1 U185 ( .Z(N1092), .A(N597) );
inv_1 U186 ( .Z(N1104), .A(N598) );
inv_1 U187 ( .Z(N1137), .A(N545) );
inv_1 U188 ( .Z(N1138), .A(N348) );
inv_1 U189 ( .Z(N1139), .A(N366) );
and2_1 U190 ( .Z(N1140), .A(N552), .B(N562) );
inv_1 U191 ( .Z(N1141), .A(N549) );
inv_1 U192 ( .Z(N1142), .A(N545) );
inv_1 U193 ( .Z(N1143), .A(N545) );
inv_1 U194 ( .Z(N1144), .A(N338) );
inv_1 U195 ( .Z(N1145), .A(N358) );
nand2_1 U196 ( .Z(N1146), .A(N373), .B(N1) );
and2_1 U197 ( .Z(N1147), .A(N141), .B(N145) );
inv_1 U198 ( .Z(N1148), .A(N592) );
inv_1 U199 ( .Z(N1149), .A(N1042) );
and2_1 U200 ( .Z(N1150), .A(N1043), .B(N27) );
and2_1 U201 ( .Z(N1151), .A(N386), .B(N556) );
inv_1 U202 ( .Z(N1152), .A(N245) );
inv_1 U203 ( .Z(N1153), .A(N552) );
inv_1 U204 ( .Z(N1154), .A(N562) );
inv_1 U205 ( .Z(N1155), .A(N559) );
and4_1 U206 ( .Z(N1156), .A(N386), .B(N559), .C(N556), .D(N552) );
inv_1 U207 ( .Z(N1157), .A(N566) );
buf_1 U208 ( .Z(N1161), .A(N571) );
buf_1 U209 ( .Z(N1173), .A(N574) );
buf_1 U210 ( .Z(N1185), .A(N571) );
buf_1 U211 ( .Z(N1197), .A(N574) );
buf_1 U212 ( .Z(N1209), .A(N137) );
buf_1 U213 ( .Z(N1213), .A(N137) );
buf_1 U214 ( .Z(N1216), .A(N141) );
inv_1 U215 ( .Z(N1219), .A(N583) );
buf_1 U216 ( .Z(N1223), .A(N577) );
buf_1 U217 ( .Z(N1235), .A(N580) );
buf_1 U218 ( .Z(N1247), .A(N577) );
buf_1 U219 ( .Z(N1259), .A(N580) );
buf_1 U220 ( .Z(N1271), .A(N254) );
buf_1 U221 ( .Z(N1280), .A(N251) );
buf_1 U222 ( .Z(N1292), .A(N251) );
buf_1 U223 ( .Z(N1303), .A(N248) );
buf_1 U224 ( .Z(N1315), .A(N248) );
buf_1 U225 ( .Z(N1327), .A(N610) );
buf_1 U226 ( .Z(N1339), .A(N607) );
buf_1 U227 ( .Z(N1351), .A(N613) );
buf_1 U228 ( .Z(N1363), .A(N616) );
buf_1 U229 ( .Z(N1375), .A(N210) );
buf_1 U230 ( .Z(N1378), .A(N210) );
buf_1 U231 ( .Z(N1381), .A(N218) );
buf_1 U232 ( .Z(N1384), .A(N218) );
buf_1 U233 ( .Z(N1387), .A(N226) );
buf_1 U234 ( .Z(N1390), .A(N226) );
buf_1 U235 ( .Z(N1393), .A(N234) );
buf_1 U236 ( .Z(N1396), .A(N234) );
buf_1 U237 ( .Z(N1415), .A(N257) );
buf_1 U238 ( .Z(N1418), .A(N257) );
buf_1 U239 ( .Z(N1421), .A(N265) );
buf_1 U240 ( .Z(N1424), .A(N265) );
buf_1 U241 ( .Z(N1427), .A(N273) );
buf_1 U242 ( .Z(N1430), .A(N273) );
buf_1 U243 ( .Z(N1433), .A(N281) );
buf_1 U244 ( .Z(N1436), .A(N281) );
buf_1 U245 ( .Z(N1455), .A(N335) );
buf_1 U246 ( .Z(N1462), .A(N335) );
buf_1 U247 ( .Z(N1469), .A(N206) );
and2_1 U248 ( .Z(N1475), .A(N27), .B(N31) );
buf_1 U249 ( .Z(N1479), .A(N1) );
buf_1 U250 ( .Z(N1482), .A(N588) );
buf_1 U251 ( .Z(N1492), .A(N293) );
buf_1 U252 ( .Z(N1495), .A(N302) );
buf_1 U253 ( .Z(N1498), .A(N308) );
buf_1 U254 ( .Z(N1501), .A(N308) );
buf_1 U255 ( .Z(N1504), .A(N316) );
buf_1 U256 ( .Z(N1507), .A(N316) );
buf_1 U257 ( .Z(N1510), .A(N324) );
buf_1 U258 ( .Z(N1513), .A(N324) );
buf_1 U259 ( .Z(N1516), .A(N341) );
buf_1 U260 ( .Z(N1519), .A(N341) );
buf_1 U261 ( .Z(N1522), .A(N351) );
buf_1 U262 ( .Z(N1525), .A(N351) );
buf_1 U263 ( .Z(N1542), .A(N257) );
buf_1 U264 ( .Z(N1545), .A(N257) );
buf_1 U265 ( .Z(N1548), .A(N265) );
buf_1 U266 ( .Z(N1551), .A(N265) );
buf_1 U267 ( .Z(N1554), .A(N273) );
buf_1 U268 ( .Z(N1557), .A(N273) );
buf_1 U269 ( .Z(N1560), .A(N281) );
buf_1 U270 ( .Z(N1563), .A(N281) );
buf_1 U271 ( .Z(N1566), .A(N332) );
buf_1 U272 ( .Z(N1573), .A(N332) );
buf_1 U273 ( .Z(N1580), .A(N549) );
and2_1 U274 ( .Z(N1583), .A(N31), .B(N27) );
inv_1 U275 ( .Z(N1588), .A(N588) );
buf_1 U276 ( .Z(N1594), .A(N324) );
buf_1 U277 ( .Z(N1597), .A(N324) );
buf_1 U278 ( .Z(N1600), .A(N341) );
buf_1 U279 ( .Z(N1603), .A(N341) );
buf_1 U280 ( .Z(N1606), .A(N351) );
buf_1 U281 ( .Z(N1609), .A(N351) );
buf_1 U282 ( .Z(N1612), .A(N293) );
buf_1 U283 ( .Z(N1615), .A(N302) );
buf_1 U284 ( .Z(N1618), .A(N308) );
buf_1 U285 ( .Z(N1621), .A(N308) );
buf_1 U286 ( .Z(N1624), .A(N316) );
buf_1 U287 ( .Z(N1627), .A(N316) );
buf_1 U288 ( .Z(N1630), .A(N361) );
buf_1 U289 ( .Z(N1633), .A(N361) );
buf_1 U290 ( .Z(N1636), .A(N210) );
buf_1 U291 ( .Z(N1639), .A(N210) );
buf_1 U292 ( .Z(N1642), .A(N218) );
buf_1 U293 ( .Z(N1645), .A(N218) );
buf_1 U294 ( .Z(N1648), .A(N226) );
buf_1 U295 ( .Z(N1651), .A(N226) );
buf_1 U296 ( .Z(N1654), .A(N234) );
buf_1 U297 ( .Z(N1657), .A(N234) );
inv_1 U298 ( .Z(N1660), .A(N324) );
buf_1 U299 ( .Z(N1663), .A(N242) );
buf_1 U300 ( .Z(N1675), .A(N242) );
buf_1 U301 ( .Z(N1685), .A(N254) );
buf_1 U302 ( .Z(N1697), .A(N610) );
buf_1 U303 ( .Z(N1709), .A(N607) );
buf_1 U304 ( .Z(N1721), .A(N625) );
buf_1 U305 ( .Z(N1727), .A(N619) );
buf_1 U306 ( .Z(N1731), .A(N613) );
buf_1 U307 ( .Z(N1743), .A(N616) );
inv_1 U308 ( .Z(N1755), .A(N599) );
inv_1 U309 ( .Z(N1758), .A(N603) );
buf_1 U310 ( .Z(N1761), .A(N619) );
buf_1 U311 ( .Z(N1769), .A(N625) );
buf_1 U312 ( .Z(N1777), .A(N619) );
buf_1 U313 ( .Z(N1785), .A(N625) );
buf_1 U314 ( .Z(N1793), .A(N619) );
buf_1 U315 ( .Z(N1800), .A(N625) );
buf_1 U316 ( .Z(N1807), .A(N619) );
buf_1 U317 ( .Z(N1814), .A(N625) );
buf_1 U318 ( .Z(N1821), .A(N299) );
buf_1 U319 ( .Z(N1824), .A(N446) );
buf_1 U320 ( .Z(N1827), .A(N457) );
buf_1 U321 ( .Z(N1830), .A(N468) );
buf_1 U322 ( .Z(N1833), .A(N422) );
buf_1 U323 ( .Z(N1836), .A(N435) );
buf_1 U324 ( .Z(N1839), .A(N389) );
buf_1 U325 ( .Z(N1842), .A(N400) );
buf_1 U326 ( .Z(N1845), .A(N411) );
buf_1 U327 ( .Z(N1848), .A(N374) );
buf_1 U328 ( .Z(N1851), .A(N4) );
buf_1 U329 ( .Z(N1854), .A(N446) );
buf_1 U330 ( .Z(N1857), .A(N457) );
buf_1 U331 ( .Z(N1860), .A(N468) );
buf_1 U332 ( .Z(N1863), .A(N435) );
buf_1 U333 ( .Z(N1866), .A(N389) );
buf_1 U334 ( .Z(N1869), .A(N400) );
buf_1 U335 ( .Z(N1872), .A(N411) );
buf_1 U336 ( .Z(N1875), .A(N422) );
buf_1 U337 ( .Z(N1878), .A(N374) );
buf_1 U338 ( .Z(N1881), .A(N479) );
buf_1 U339 ( .Z(N1884), .A(N490) );
buf_1 U340 ( .Z(N1887), .A(N503) );
buf_1 U341 ( .Z(N1890), .A(N514) );
buf_1 U342 ( .Z(N1893), .A(N523) );
buf_1 U343 ( .Z(N1896), .A(N534) );
buf_1 U344 ( .Z(N1899), .A(N54) );
buf_1 U345 ( .Z(N1902), .A(N479) );
buf_1 U346 ( .Z(N1905), .A(N503) );
buf_1 U347 ( .Z(N1908), .A(N514) );
buf_1 U348 ( .Z(N1911), .A(N523) );
buf_1 U349 ( .Z(N1914), .A(N534) );
buf_1 U350 ( .Z(N1917), .A(N490) );
buf_1 U351 ( .Z(N1920), .A(N361) );
buf_1 U352 ( .Z(N1923), .A(N369) );
buf_1 U353 ( .Z(N1926), .A(N341) );
buf_1 U354 ( .Z(N1929), .A(N351) );
buf_1 U355 ( .Z(N1932), .A(N308) );
buf_1 U356 ( .Z(N1935), .A(N316) );
buf_1 U357 ( .Z(N1938), .A(N293) );
buf_1 U358 ( .Z(N1941), .A(N302) );
buf_1 U359 ( .Z(N1944), .A(N281) );
buf_1 U360 ( .Z(N1947), .A(N289) );
buf_1 U361 ( .Z(N1950), .A(N265) );
buf_1 U362 ( .Z(N1953), .A(N273) );
buf_1 U363 ( .Z(N1956), .A(N234) );
buf_1 U364 ( .Z(N1959), .A(N257) );
buf_1 U365 ( .Z(N1962), .A(N218) );
buf_1 U366 ( .Z(N1965), .A(N226) );
buf_1 U367 ( .Z(N1968), .A(N210) );
inv_1 U368 ( .Z(N1972), .A(N1146) );
and2_1 U369 ( .Z(N2054), .A(N136), .B(N1148) );
inv_1 U370 ( .Z(N2060), .A(N1150) );
inv_1 U371 ( .Z(N2061), .A(N1151) );
buf_1 U372 ( .Z(N2139), .A(N1209) );
buf_1 U373 ( .Z(N2142), .A(N1216) );
buf_1 U374 ( .Z(N2309), .A(N1479) );
and2_1 U375 ( .Z(N2349), .A(N1104), .B(N514) );
or2_1 U376 ( .Z(N2350), .A(N1067), .B(N514) );
buf_1 U377 ( .Z(N2387), .A(N1580) );
buf_1 U378 ( .Z(N2527), .A(N1821) );
inv_1 U379 ( .Z(N2584), .A(N1580) );
and3_1 U380 ( .Z(N2585), .A(N170), .B(N1161), .C(N1173) );
and3_1 U381 ( .Z(N2586), .A(N173), .B(N1161), .C(N1173) );
and3_1 U382 ( .Z(N2587), .A(N167), .B(N1161), .C(N1173) );
and3_1 U383 ( .Z(N2588), .A(N164), .B(N1161), .C(N1173) );
and3_1 U384 ( .Z(N2589), .A(N161), .B(N1161), .C(N1173) );
nand2_1 U385 ( .Z(N2590), .A(N1475), .B(N140) );
and3_1 U386 ( .Z(N2591), .A(N185), .B(N1185), .C(N1197) );
and3_1 U387 ( .Z(N2592), .A(N158), .B(N1185), .C(N1197) );
and3_1 U388 ( .Z(N2593), .A(N152), .B(N1185), .C(N1197) );
and3_1 U389 ( .Z(N2594), .A(N146), .B(N1185), .C(N1197) );
and3_1 U390 ( .Z(N2595), .A(N170), .B(N1223), .C(N1235) );
and3_1 U391 ( .Z(N2596), .A(N173), .B(N1223), .C(N1235) );
and3_1 U392 ( .Z(N2597), .A(N167), .B(N1223), .C(N1235) );
and3_1 U393 ( .Z(N2598), .A(N164), .B(N1223), .C(N1235) );
and3_1 U394 ( .Z(N2599), .A(N161), .B(N1223), .C(N1235) );
and3_1 U395 ( .Z(N2600), .A(N185), .B(N1247), .C(N1259) );
and3_1 U396 ( .Z(N2601), .A(N158), .B(N1247), .C(N1259) );
and3_1 U397 ( .Z(N2602), .A(N152), .B(N1247), .C(N1259) );
and3_1 U398 ( .Z(N2603), .A(N146), .B(N1247), .C(N1259) );
and3_1 U399 ( .Z(N2604), .A(N106), .B(N1731), .C(N1743) );
and3_1 U400 ( .Z(N2605), .A(N61), .B(N1327), .C(N1339) );
and3_1 U401 ( .Z(N2606), .A(N106), .B(N1697), .C(N1709) );
and3_1 U402 ( .Z(N2607), .A(N49), .B(N1697), .C(N1709) );
and3_1 U403 ( .Z(N2608), .A(N103), .B(N1697), .C(N1709) );
and3_1 U404 ( .Z(N2609), .A(N40), .B(N1697), .C(N1709) );
and3_1 U405 ( .Z(N2610), .A(N37), .B(N1697), .C(N1709) );
and3_1 U406 ( .Z(N2611), .A(N20), .B(N1327), .C(N1339) );
and3_1 U407 ( .Z(N2612), .A(N17), .B(N1327), .C(N1339) );
and3_1 U408 ( .Z(N2613), .A(N70), .B(N1327), .C(N1339) );
and3_1 U409 ( .Z(N2614), .A(N64), .B(N1327), .C(N1339) );
and3_1 U410 ( .Z(N2615), .A(N49), .B(N1731), .C(N1743) );
and3_1 U411 ( .Z(N2616), .A(N103), .B(N1731), .C(N1743) );
and3_1 U412 ( .Z(N2617), .A(N40), .B(N1731), .C(N1743) );
and3_1 U413 ( .Z(N2618), .A(N37), .B(N1731), .C(N1743) );
and3_1 U414 ( .Z(N2619), .A(N20), .B(N1351), .C(N1363) );
and3_1 U415 ( .Z(N2620), .A(N17), .B(N1351), .C(N1363) );
and3_1 U416 ( .Z(N2621), .A(N70), .B(N1351), .C(N1363) );
and3_1 U417 ( .Z(N2622), .A(N64), .B(N1351), .C(N1363) );
inv_1 U418 ( .Z(N2623), .A(N1475) );
and3_1 U419 ( .Z(N2624), .A(N123), .B(N1758), .C(N599) );
and2_1 U420 ( .Z(N2625), .A(N1777), .B(N1785) );
and3_1 U421 ( .Z(N2626), .A(N61), .B(N1351), .C(N1363) );
and2_1 U422 ( .Z(N2627), .A(N1761), .B(N1769) );
inv_1 U423 ( .Z(N2628), .A(N1824) );
inv_1 U424 ( .Z(N2629), .A(N1827) );
inv_1 U425 ( .Z(N2630), .A(N1830) );
inv_1 U426 ( .Z(N2631), .A(N1833) );
inv_1 U427 ( .Z(N2632), .A(N1836) );
inv_1 U428 ( .Z(N2633), .A(N1839) );
inv_1 U429 ( .Z(N2634), .A(N1842) );
inv_1 U430 ( .Z(N2635), .A(N1845) );
inv_1 U431 ( .Z(N2636), .A(N1848) );
inv_1 U432 ( .Z(N2637), .A(N1851) );
inv_1 U433 ( .Z(N2638), .A(N1854) );
inv_1 U434 ( .Z(N2639), .A(N1857) );
inv_1 U435 ( .Z(N2640), .A(N1860) );
inv_1 U436 ( .Z(N2641), .A(N1863) );
inv_1 U437 ( .Z(N2642), .A(N1866) );
inv_1 U438 ( .Z(N2643), .A(N1869) );
inv_1 U439 ( .Z(N2644), .A(N1872) );
inv_1 U440 ( .Z(N2645), .A(N1875) );
inv_1 U441 ( .Z(N2646), .A(N1878) );
buf_1 U442 ( .Z(N2647), .A(N1209) );
inv_1 U443 ( .Z(N2653), .A(N1161) );
inv_1 U444 ( .Z(N2664), .A(N1173) );
buf_1 U445 ( .Z(N2675), .A(N1209) );
inv_1 U446 ( .Z(N2681), .A(N1185) );
inv_1 U447 ( .Z(N2692), .A(N1197) );
and3_1 U448 ( .Z(N2703), .A(N179), .B(N1185), .C(N1197) );
buf_1 U449 ( .Z(N2704), .A(N1479) );
inv_1 U450 ( .Z(N2709), .A(N1881) );
inv_1 U451 ( .Z(N2710), .A(N1884) );
inv_1 U452 ( .Z(N2711), .A(N1887) );
inv_1 U453 ( .Z(N2712), .A(N1890) );
inv_1 U454 ( .Z(N2713), .A(N1893) );
inv_1 U455 ( .Z(N2714), .A(N1896) );
inv_1 U456 ( .Z(N2715), .A(N1899) );
inv_1 U457 ( .Z(N2716), .A(N1902) );
inv_1 U458 ( .Z(N2717), .A(N1905) );
inv_1 U459 ( .Z(N2718), .A(N1908) );
inv_1 U460 ( .Z(N2719), .A(N1911) );
inv_1 U461 ( .Z(N2720), .A(N1914) );
inv_1 U462 ( .Z(N2721), .A(N1917) );
buf_1 U463 ( .Z(N2722), .A(N1213) );
inv_1 U464 ( .Z(N2728), .A(N1223) );
inv_1 U465 ( .Z(N2739), .A(N1235) );
buf_1 U466 ( .Z(N2750), .A(N1213) );
inv_1 U467 ( .Z(N2756), .A(N1247) );
inv_1 U468 ( .Z(N2767), .A(N1259) );
and3_1 U469 ( .Z(N2778), .A(N179), .B(N1247), .C(N1259) );
inv_1 U470 ( .Z(N2779), .A(N1327) );
inv_1 U471 ( .Z(N2790), .A(N1339) );
inv_1 U472 ( .Z(N2801), .A(N1351) );
inv_1 U473 ( .Z(N2812), .A(N1363) );
inv_1 U474 ( .Z(N2823), .A(N1375) );
inv_1 U475 ( .Z(N2824), .A(N1378) );
inv_1 U476 ( .Z(N2825), .A(N1381) );
inv_1 U477 ( .Z(N2826), .A(N1384) );
inv_1 U478 ( .Z(N2827), .A(N1387) );
inv_1 U479 ( .Z(N2828), .A(N1390) );
inv_1 U480 ( .Z(N2829), .A(N1393) );
inv_1 U481 ( .Z(N2830), .A(N1396) );
and3_1 U482 ( .Z(N2831), .A(N1104), .B(N457), .C(N1378) );
and3_1 U483 ( .Z(N2832), .A(N1104), .B(N468), .C(N1384) );
and3_1 U484 ( .Z(N2833), .A(N1104), .B(N422), .C(N1390) );
and3_1 U485 ( .Z(N2834), .A(N1104), .B(N435), .C(N1396) );
and2_1 U486 ( .Z(N2835), .A(N1067), .B(N1375) );
and2_1 U487 ( .Z(N2836), .A(N1067), .B(N1381) );
and2_1 U488 ( .Z(N2837), .A(N1067), .B(N1387) );
and2_1 U489 ( .Z(N2838), .A(N1067), .B(N1393) );
inv_1 U490 ( .Z(N2839), .A(N1415) );
inv_1 U491 ( .Z(N2840), .A(N1418) );
inv_1 U492 ( .Z(N2841), .A(N1421) );
inv_1 U493 ( .Z(N2842), .A(N1424) );
inv_1 U494 ( .Z(N2843), .A(N1427) );
inv_1 U495 ( .Z(N2844), .A(N1430) );
inv_1 U496 ( .Z(N2845), .A(N1433) );
inv_1 U497 ( .Z(N2846), .A(N1436) );
and3_1 U498 ( .Z(N2847), .A(N1104), .B(N389), .C(N1418) );
and3_1 U499 ( .Z(N2848), .A(N1104), .B(N400), .C(N1424) );
and3_1 U500 ( .Z(N2849), .A(N1104), .B(N411), .C(N1430) );
and3_1 U501 ( .Z(N2850), .A(N1104), .B(N374), .C(N1436) );
and2_1 U502 ( .Z(N2851), .A(N1067), .B(N1415) );
and2_1 U503 ( .Z(N2852), .A(N1067), .B(N1421) );
and2_1 U504 ( .Z(N2853), .A(N1067), .B(N1427) );
and2_1 U505 ( .Z(N2854), .A(N1067), .B(N1433) );
inv_1 U506 ( .Z(N2855), .A(N1455) );
inv_1 U507 ( .Z(N2861), .A(N1462) );
and2_1 U508 ( .Z(N2867), .A(N292), .B(N1455) );
and2_1 U509 ( .Z(N2868), .A(N288), .B(N1455) );
and2_1 U510 ( .Z(N2869), .A(N280), .B(N1455) );
and2_1 U511 ( .Z(N2870), .A(N272), .B(N1455) );
and2_1 U512 ( .Z(N2871), .A(N264), .B(N1455) );
and2_1 U513 ( .Z(N2872), .A(N241), .B(N1462) );
and2_1 U514 ( .Z(N2873), .A(N233), .B(N1462) );
and2_1 U515 ( .Z(N2874), .A(N225), .B(N1462) );
and2_1 U516 ( .Z(N2875), .A(N217), .B(N1462) );
and2_1 U517 ( .Z(N2876), .A(N209), .B(N1462) );
buf_1 U518 ( .Z(N2877), .A(N1216) );
inv_1 U519 ( .Z(N2882), .A(N1482) );
inv_1 U520 ( .Z(N2891), .A(N1475) );
inv_1 U521 ( .Z(N2901), .A(N1492) );
inv_1 U522 ( .Z(N2902), .A(N1495) );
inv_1 U523 ( .Z(N2903), .A(N1498) );
inv_1 U524 ( .Z(N2904), .A(N1501) );
inv_1 U525 ( .Z(N2905), .A(N1504) );
inv_1 U526 ( .Z(N2906), .A(N1507) );
and2_1 U527 ( .Z(N2907), .A(N1303), .B(N1495) );
and3_1 U528 ( .Z(N2908), .A(N1303), .B(N479), .C(N1501) );
and3_1 U529 ( .Z(N2909), .A(N1303), .B(N490), .C(N1507) );
and2_1 U530 ( .Z(N2910), .A(N1663), .B(N1492) );
and2_1 U531 ( .Z(N2911), .A(N1663), .B(N1498) );
and2_1 U532 ( .Z(N2912), .A(N1663), .B(N1504) );
inv_1 U533 ( .Z(N2913), .A(N1510) );
inv_1 U534 ( .Z(N2914), .A(N1513) );
inv_1 U535 ( .Z(N2915), .A(N1516) );
inv_1 U536 ( .Z(N2916), .A(N1519) );
inv_1 U537 ( .Z(N2917), .A(N1522) );
inv_1 U538 ( .Z(N2918), .A(N1525) );
and3_1 U539 ( .Z(N2919), .A(N1104), .B(N503), .C(N1513) );
inv_1 U540 ( .Z(N2920), .A(N2349) );
and3_1 U541 ( .Z(N2921), .A(N1104), .B(N523), .C(N1519) );
and3_1 U542 ( .Z(N2922), .A(N1104), .B(N534), .C(N1525) );
and2_1 U543 ( .Z(N2923), .A(N1067), .B(N1510) );
and2_1 U544 ( .Z(N2924), .A(N1067), .B(N1516) );
and2_1 U545 ( .Z(N2925), .A(N1067), .B(N1522) );
inv_1 U546 ( .Z(N2926), .A(N1542) );
inv_1 U547 ( .Z(N2927), .A(N1545) );
inv_1 U548 ( .Z(N2928), .A(N1548) );
inv_1 U549 ( .Z(N2929), .A(N1551) );
inv_1 U550 ( .Z(N2930), .A(N1554) );
inv_1 U551 ( .Z(N2931), .A(N1557) );
inv_1 U552 ( .Z(N2932), .A(N1560) );
inv_1 U553 ( .Z(N2933), .A(N1563) );
and3_1 U554 ( .Z(N2934), .A(N1303), .B(N389), .C(N1545) );
and3_1 U555 ( .Z(N2935), .A(N1303), .B(N400), .C(N1551) );
and3_1 U556 ( .Z(N2936), .A(N1303), .B(N411), .C(N1557) );
and3_1 U557 ( .Z(N2937), .A(N1303), .B(N374), .C(N1563) );
and2_1 U558 ( .Z(N2938), .A(N1663), .B(N1542) );
and2_1 U559 ( .Z(N2939), .A(N1663), .B(N1548) );
and2_1 U560 ( .Z(N2940), .A(N1663), .B(N1554) );
and2_1 U561 ( .Z(N2941), .A(N1663), .B(N1560) );
inv_1 U562 ( .Z(N2942), .A(N1566) );
inv_1 U563 ( .Z(N2948), .A(N1573) );
and2_1 U564 ( .Z(N2954), .A(N372), .B(N1566) );
and2_1 U565 ( .Z(N2955), .A(N366), .B(N1566) );
and2_1 U566 ( .Z(N2956), .A(N358), .B(N1566) );
and2_1 U567 ( .Z(N2957), .A(N348), .B(N1566) );
and2_1 U568 ( .Z(N2958), .A(N338), .B(N1566) );
and2_1 U569 ( .Z(N2959), .A(N331), .B(N1573) );
and2_1 U570 ( .Z(N2960), .A(N323), .B(N1573) );
and2_1 U571 ( .Z(N2961), .A(N315), .B(N1573) );
and2_1 U572 ( .Z(N2962), .A(N307), .B(N1573) );
and2_1 U573 ( .Z(N2963), .A(N299), .B(N1573) );
inv_1 U574 ( .Z(N2964), .A(N1588) );
and2_1 U575 ( .Z(N2969), .A(N83), .B(N1588) );
and2_1 U576 ( .Z(N2970), .A(N86), .B(N1588) );
and2_1 U577 ( .Z(N2971), .A(N88), .B(N1588) );
and2_1 U578 ( .Z(N2972), .A(N88), .B(N1588) );
inv_1 U579 ( .Z(N2973), .A(N1594) );
inv_1 U580 ( .Z(N2974), .A(N1597) );
inv_1 U581 ( .Z(N2975), .A(N1600) );
inv_1 U582 ( .Z(N2976), .A(N1603) );
inv_1 U583 ( .Z(N2977), .A(N1606) );
inv_1 U584 ( .Z(N2978), .A(N1609) );
and3_1 U585 ( .Z(N2979), .A(N1315), .B(N503), .C(N1597) );
and2_1 U586 ( .Z(N2980), .A(N1315), .B(N514) );
and3_1 U587 ( .Z(N2981), .A(N1315), .B(N523), .C(N1603) );
and3_1 U588 ( .Z(N2982), .A(N1315), .B(N534), .C(N1609) );
and2_1 U589 ( .Z(N2983), .A(N1675), .B(N1594) );
or2_1 U590 ( .Z(N2984), .A(N1675), .B(N514) );
and2_1 U591 ( .Z(N2985), .A(N1675), .B(N1600) );
and2_1 U592 ( .Z(N2986), .A(N1675), .B(N1606) );
inv_1 U593 ( .Z(N2987), .A(N1612) );
inv_1 U594 ( .Z(N2988), .A(N1615) );
inv_1 U595 ( .Z(N2989), .A(N1618) );
inv_1 U596 ( .Z(N2990), .A(N1621) );
inv_1 U597 ( .Z(N2991), .A(N1624) );
inv_1 U598 ( .Z(N2992), .A(N1627) );
and2_1 U599 ( .Z(N2993), .A(N1315), .B(N1615) );
and3_1 U600 ( .Z(N2994), .A(N1315), .B(N479), .C(N1621) );
and3_1 U601 ( .Z(N2995), .A(N1315), .B(N490), .C(N1627) );
and2_1 U602 ( .Z(N2996), .A(N1675), .B(N1612) );
and2_1 U603 ( .Z(N2997), .A(N1675), .B(N1618) );
and2_1 U604 ( .Z(N2998), .A(N1675), .B(N1624) );
inv_1 U605 ( .Z(N2999), .A(N1630) );
buf_1 U606 ( .Z(N3000), .A(N1469) );
buf_1 U607 ( .Z(N3003), .A(N1469) );
inv_1 U608 ( .Z(N3006), .A(N1633) );
buf_1 U609 ( .Z(N3007), .A(N1469) );
buf_1 U610 ( .Z(N3010), .A(N1469) );
and2_1 U611 ( .Z(N3013), .A(N1315), .B(N1630) );
and2_1 U612 ( .Z(N3014), .A(N1315), .B(N1633) );
inv_1 U613 ( .Z(N3015), .A(N1636) );
inv_1 U614 ( .Z(N3016), .A(N1639) );
inv_1 U615 ( .Z(N3017), .A(N1642) );
inv_1 U616 ( .Z(N3018), .A(N1645) );
inv_1 U617 ( .Z(N3019), .A(N1648) );
inv_1 U618 ( .Z(N3020), .A(N1651) );
inv_1 U619 ( .Z(N3021), .A(N1654) );
inv_1 U620 ( .Z(N3022), .A(N1657) );
and3_1 U621 ( .Z(N3023), .A(N1303), .B(N457), .C(N1639) );
and3_1 U622 ( .Z(N3024), .A(N1303), .B(N468), .C(N1645) );
and3_1 U623 ( .Z(N3025), .A(N1303), .B(N422), .C(N1651) );
and3_1 U624 ( .Z(N3026), .A(N1303), .B(N435), .C(N1657) );
and2_1 U625 ( .Z(N3027), .A(N1663), .B(N1636) );
and2_1 U626 ( .Z(N3028), .A(N1663), .B(N1642) );
and2_1 U627 ( .Z(N3029), .A(N1663), .B(N1648) );
and2_1 U628 ( .Z(N3030), .A(N1663), .B(N1654) );
inv_1 U629 ( .Z(N3031), .A(N1920) );
inv_1 U630 ( .Z(N3032), .A(N1923) );
inv_1 U631 ( .Z(N3033), .A(N1926) );
inv_1 U632 ( .Z(N3034), .A(N1929) );
buf_1 U633 ( .Z(N3035), .A(N1660) );
buf_1 U634 ( .Z(N3038), .A(N1660) );
inv_1 U635 ( .Z(N3041), .A(N1697) );
inv_1 U636 ( .Z(N3052), .A(N1709) );
inv_1 U637 ( .Z(N3063), .A(N1721) );
inv_1 U638 ( .Z(N3068), .A(N1727) );
and2_1 U639 ( .Z(N3071), .A(N97), .B(N1721) );
and2_1 U640 ( .Z(N3072), .A(N94), .B(N1721) );
and2_1 U641 ( .Z(N3073), .A(N97), .B(N1721) );
and2_1 U642 ( .Z(N3074), .A(N94), .B(N1721) );
inv_1 U643 ( .Z(N3075), .A(N1731) );
inv_1 U644 ( .Z(N3086), .A(N1743) );
inv_1 U645 ( .Z(N3097), .A(N1761) );
inv_1 U646 ( .Z(N3108), .A(N1769) );
inv_1 U647 ( .Z(N3119), .A(N1777) );
inv_1 U648 ( .Z(N3130), .A(N1785) );
inv_1 U649 ( .Z(N3141), .A(N1944) );
inv_1 U650 ( .Z(N3142), .A(N1947) );
inv_1 U651 ( .Z(N3143), .A(N1950) );
inv_1 U652 ( .Z(N3144), .A(N1953) );
inv_1 U653 ( .Z(N3145), .A(N1956) );
inv_1 U654 ( .Z(N3146), .A(N1959) );
inv_1 U655 ( .Z(N3147), .A(N1793) );
inv_1 U656 ( .Z(N3158), .A(N1800) );
inv_1 U657 ( .Z(N3169), .A(N1807) );
inv_1 U658 ( .Z(N3180), .A(N1814) );
buf_1 U659 ( .Z(N3191), .A(N1821) );
inv_1 U660 ( .Z(N3194), .A(N1932) );
inv_1 U661 ( .Z(N3195), .A(N1935) );
inv_1 U662 ( .Z(N3196), .A(N1938) );
inv_1 U663 ( .Z(N3197), .A(N1941) );
inv_1 U664 ( .Z(N3198), .A(N1962) );
inv_1 U665 ( .Z(N3199), .A(N1965) );
buf_1 U666 ( .Z(N3200), .A(N1469) );
inv_1 U667 ( .Z(N3203), .A(N1968) );
buf_1 U668 ( .Z(N3357), .A(N2704) );
buf_1 U669 ( .Z(N3358), .A(N2704) );
buf_1 U670 ( .Z(N3359), .A(N2704) );
buf_1 U671 ( .Z(N3360), .A(N2704) );
and3_1 U672 ( .Z(N3401), .A(N457), .B(N1092), .C(N2824) );
and3_1 U673 ( .Z(N3402), .A(N468), .B(N1092), .C(N2826) );
and3_1 U674 ( .Z(N3403), .A(N422), .B(N1092), .C(N2828) );
and3_1 U675 ( .Z(N3404), .A(N435), .B(N1092), .C(N2830) );
and2_1 U676 ( .Z(N3405), .A(N1080), .B(N2823) );
and2_1 U677 ( .Z(N3406), .A(N1080), .B(N2825) );
and2_1 U678 ( .Z(N3407), .A(N1080), .B(N2827) );
and2_1 U679 ( .Z(N3408), .A(N1080), .B(N2829) );
and3_1 U680 ( .Z(N3409), .A(N389), .B(N1092), .C(N2840) );
and3_1 U681 ( .Z(N3410), .A(N400), .B(N1092), .C(N2842) );
and3_1 U682 ( .Z(N3411), .A(N411), .B(N1092), .C(N2844) );
and3_1 U683 ( .Z(N3412), .A(N374), .B(N1092), .C(N2846) );
and2_1 U684 ( .Z(N3413), .A(N1080), .B(N2839) );
and2_1 U685 ( .Z(N3414), .A(N1080), .B(N2841) );
and2_1 U686 ( .Z(N3415), .A(N1080), .B(N2843) );
and2_1 U687 ( .Z(N3416), .A(N1080), .B(N2845) );
and2_1 U688 ( .Z(N3444), .A(N1280), .B(N2902) );
and3_1 U689 ( .Z(N3445), .A(N479), .B(N1280), .C(N2904) );
and3_1 U690 ( .Z(N3446), .A(N490), .B(N1280), .C(N2906) );
and2_1 U691 ( .Z(N3447), .A(N1685), .B(N2901) );
and2_1 U692 ( .Z(N3448), .A(N1685), .B(N2903) );
and2_1 U693 ( .Z(N3449), .A(N1685), .B(N2905) );
and3_1 U694 ( .Z(N3450), .A(N503), .B(N1092), .C(N2914) );
and3_1 U695 ( .Z(N3451), .A(N523), .B(N1092), .C(N2916) );
and3_1 U696 ( .Z(N3452), .A(N534), .B(N1092), .C(N2918) );
and2_1 U697 ( .Z(N3453), .A(N1080), .B(N2913) );
and2_1 U698 ( .Z(N3454), .A(N1080), .B(N2915) );
and2_1 U699 ( .Z(N3455), .A(N1080), .B(N2917) );
and2_1 U700 ( .Z(N3456), .A(N2920), .B(N2350) );
and3_1 U701 ( .Z(N3459), .A(N389), .B(N1280), .C(N2927) );
and3_1 U702 ( .Z(N3460), .A(N400), .B(N1280), .C(N2929) );
and3_1 U703 ( .Z(N3461), .A(N411), .B(N1280), .C(N2931) );
and3_1 U704 ( .Z(N3462), .A(N374), .B(N1280), .C(N2933) );
and2_1 U705 ( .Z(N3463), .A(N1685), .B(N2926) );
and2_1 U706 ( .Z(N3464), .A(N1685), .B(N2928) );
and2_1 U707 ( .Z(N3465), .A(N1685), .B(N2930) );
and2_1 U708 ( .Z(N3466), .A(N1685), .B(N2932) );
and3_1 U709 ( .Z(N3481), .A(N503), .B(N1292), .C(N2974) );
inv_1 U710 ( .Z(N3482), .A(N2980) );
and3_1 U711 ( .Z(N3483), .A(N523), .B(N1292), .C(N2976) );
and3_1 U712 ( .Z(N3484), .A(N534), .B(N1292), .C(N2978) );
and2_1 U713 ( .Z(N3485), .A(N1271), .B(N2973) );
and2_1 U714 ( .Z(N3486), .A(N1271), .B(N2975) );
and2_1 U715 ( .Z(N3487), .A(N1271), .B(N2977) );
and2_1 U716 ( .Z(N3488), .A(N1292), .B(N2988) );
and3_1 U717 ( .Z(N3489), .A(N479), .B(N1292), .C(N2990) );
and3_1 U718 ( .Z(N3490), .A(N490), .B(N1292), .C(N2992) );
and2_1 U719 ( .Z(N3491), .A(N1271), .B(N2987) );
and2_1 U720 ( .Z(N3492), .A(N1271), .B(N2989) );
and2_1 U721 ( .Z(N3493), .A(N1271), .B(N2991) );
and2_1 U722 ( .Z(N3502), .A(N1292), .B(N2999) );
and2_1 U723 ( .Z(N3503), .A(N1292), .B(N3006) );
and3_1 U724 ( .Z(N3504), .A(N457), .B(N1280), .C(N3016) );
and3_1 U725 ( .Z(N3505), .A(N468), .B(N1280), .C(N3018) );
and3_1 U726 ( .Z(N3506), .A(N422), .B(N1280), .C(N3020) );
and3_1 U727 ( .Z(N3507), .A(N435), .B(N1280), .C(N3022) );
and2_1 U728 ( .Z(N3508), .A(N1685), .B(N3015) );
and2_1 U729 ( .Z(N3509), .A(N1685), .B(N3017) );
and2_1 U730 ( .Z(N3510), .A(N1685), .B(N3019) );
and2_1 U731 ( .Z(N3511), .A(N1685), .B(N3021) );
nand2_1 U732 ( .Z(N3512), .A(N1923), .B(N3031) );
nand2_1 U733 ( .Z(N3513), .A(N1920), .B(N3032) );
nand2_1 U734 ( .Z(N3514), .A(N1929), .B(N3033) );
nand2_1 U735 ( .Z(N3515), .A(N1926), .B(N3034) );
nand2_1 U736 ( .Z(N3558), .A(N1947), .B(N3141) );
nand2_1 U737 ( .Z(N3559), .A(N1944), .B(N3142) );
nand2_1 U738 ( .Z(N3560), .A(N1953), .B(N3143) );
nand2_1 U739 ( .Z(N3561), .A(N1950), .B(N3144) );
nand2_1 U740 ( .Z(N3562), .A(N1959), .B(N3145) );
nand2_1 U741 ( .Z(N3563), .A(N1956), .B(N3146) );
buf_1 U742 ( .Z(N3604), .A(N3191) );
nand2_1 U743 ( .Z(N3605), .A(N1935), .B(N3194) );
nand2_1 U744 ( .Z(N3606), .A(N1932), .B(N3195) );
nand2_1 U745 ( .Z(N3607), .A(N1941), .B(N3196) );
nand2_1 U746 ( .Z(N3608), .A(N1938), .B(N3197) );
nand2_1 U747 ( .Z(N3609), .A(N1965), .B(N3198) );
nand2_1 U748 ( .Z(N3610), .A(N1962), .B(N3199) );
inv_1 U749 ( .Z(N3613), .A(N3191) );
and2_1 U750 ( .Z(N3614), .A(N2882), .B(N2891) );
and2_1 U751 ( .Z(N3615), .A(N1482), .B(N2891) );
and3_1 U752 ( .Z(N3616), .A(N200), .B(N2653), .C(N1173) );
and3_1 U753 ( .Z(N3617), .A(N203), .B(N2653), .C(N1173) );
and3_1 U754 ( .Z(N3618), .A(N197), .B(N2653), .C(N1173) );
and3_1 U755 ( .Z(N3619), .A(N194), .B(N2653), .C(N1173) );
and3_1 U756 ( .Z(N3620), .A(N191), .B(N2653), .C(N1173) );
and3_1 U757 ( .Z(N3621), .A(N182), .B(N2681), .C(N1197) );
and3_1 U758 ( .Z(N3622), .A(N188), .B(N2681), .C(N1197) );
and3_1 U759 ( .Z(N3623), .A(N155), .B(N2681), .C(N1197) );
and3_1 U760 ( .Z(N3624), .A(N149), .B(N2681), .C(N1197) );
and2_1 U761 ( .Z(N3625), .A(N2882), .B(N2891) );
and2_1 U762 ( .Z(N3626), .A(N1482), .B(N2891) );
and3_1 U763 ( .Z(N3627), .A(N200), .B(N2728), .C(N1235) );
and3_1 U764 ( .Z(N3628), .A(N203), .B(N2728), .C(N1235) );
and3_1 U765 ( .Z(N3629), .A(N197), .B(N2728), .C(N1235) );
and3_1 U766 ( .Z(N3630), .A(N194), .B(N2728), .C(N1235) );
and3_1 U767 ( .Z(N3631), .A(N191), .B(N2728), .C(N1235) );
and3_1 U768 ( .Z(N3632), .A(N182), .B(N2756), .C(N1259) );
and3_1 U769 ( .Z(N3633), .A(N188), .B(N2756), .C(N1259) );
and3_1 U770 ( .Z(N3634), .A(N155), .B(N2756), .C(N1259) );
and3_1 U771 ( .Z(N3635), .A(N149), .B(N2756), .C(N1259) );
and2_1 U772 ( .Z(N3636), .A(N2882), .B(N2891) );
and2_1 U773 ( .Z(N3637), .A(N1482), .B(N2891) );
and3_1 U774 ( .Z(N3638), .A(N109), .B(N3075), .C(N1743) );
and2_1 U775 ( .Z(N3639), .A(N2882), .B(N2891) );
and2_1 U776 ( .Z(N3640), .A(N1482), .B(N2891) );
and3_1 U777 ( .Z(N3641), .A(N11), .B(N2779), .C(N1339) );
and3_1 U778 ( .Z(N3642), .A(N109), .B(N3041), .C(N1709) );
and3_1 U779 ( .Z(N3643), .A(N46), .B(N3041), .C(N1709) );
and3_1 U780 ( .Z(N3644), .A(N100), .B(N3041), .C(N1709) );
and3_1 U781 ( .Z(N3645), .A(N91), .B(N3041), .C(N1709) );
and3_1 U782 ( .Z(N3646), .A(N43), .B(N3041), .C(N1709) );
and3_1 U783 ( .Z(N3647), .A(N76), .B(N2779), .C(N1339) );
and3_1 U784 ( .Z(N3648), .A(N73), .B(N2779), .C(N1339) );
and3_1 U785 ( .Z(N3649), .A(N67), .B(N2779), .C(N1339) );
and3_1 U786 ( .Z(N3650), .A(N14), .B(N2779), .C(N1339) );
and3_1 U787 ( .Z(N3651), .A(N46), .B(N3075), .C(N1743) );
and3_1 U788 ( .Z(N3652), .A(N100), .B(N3075), .C(N1743) );
and3_1 U789 ( .Z(N3653), .A(N91), .B(N3075), .C(N1743) );
and3_1 U790 ( .Z(N3654), .A(N43), .B(N3075), .C(N1743) );
and3_1 U791 ( .Z(N3655), .A(N76), .B(N2801), .C(N1363) );
and3_1 U792 ( .Z(N3656), .A(N73), .B(N2801), .C(N1363) );
and3_1 U793 ( .Z(N3657), .A(N67), .B(N2801), .C(N1363) );
and3_1 U794 ( .Z(N3658), .A(N14), .B(N2801), .C(N1363) );
and3_1 U795 ( .Z(N3659), .A(N120), .B(N3119), .C(N1785) );
and3_1 U796 ( .Z(N3660), .A(N11), .B(N2801), .C(N1363) );
and3_1 U797 ( .Z(N3661), .A(N118), .B(N3097), .C(N1769) );
and3_1 U798 ( .Z(N3662), .A(N176), .B(N2681), .C(N1197) );
and3_1 U799 ( .Z(N3663), .A(N176), .B(N2756), .C(N1259) );
or2_1 U800 ( .Z(N3664), .A(N2831), .B(N3401) );
or2_1 U801 ( .Z(N3665), .A(N2832), .B(N3402) );
or2_1 U802 ( .Z(N3666), .A(N2833), .B(N3403) );
or2_1 U803 ( .Z(N3667), .A(N2834), .B(N3404) );
or3_1 U804 ( .Z(N3668), .A(N2835), .B(N3405), .C(N457) );
or3_1 U805 ( .Z(N3669), .A(N2836), .B(N3406), .C(N468) );
or3_1 U806 ( .Z(N3670), .A(N2837), .B(N3407), .C(N422) );
or3_1 U807 ( .Z(N3671), .A(N2838), .B(N3408), .C(N435) );
or2_1 U808 ( .Z(N3672), .A(N2847), .B(N3409) );
or2_1 U809 ( .Z(N3673), .A(N2848), .B(N3410) );
or2_1 U810 ( .Z(N3674), .A(N2849), .B(N3411) );
or2_1 U811 ( .Z(N3675), .A(N2850), .B(N3412) );
or3_1 U812 ( .Z(N3676), .A(N2851), .B(N3413), .C(N389) );
or3_1 U813 ( .Z(N3677), .A(N2852), .B(N3414), .C(N400) );
or3_1 U814 ( .Z(N3678), .A(N2853), .B(N3415), .C(N411) );
or3_1 U815 ( .Z(N3679), .A(N2854), .B(N3416), .C(N374) );
and2_1 U816 ( .Z(N3680), .A(N289), .B(N2855) );
and2_1 U817 ( .Z(N3681), .A(N281), .B(N2855) );
and2_1 U818 ( .Z(N3682), .A(N273), .B(N2855) );
and2_1 U819 ( .Z(N3683), .A(N265), .B(N2855) );
and2_1 U820 ( .Z(N3684), .A(N257), .B(N2855) );
and2_1 U821 ( .Z(N3685), .A(N234), .B(N2861) );
and2_1 U822 ( .Z(N3686), .A(N226), .B(N2861) );
and2_1 U823 ( .Z(N3687), .A(N218), .B(N2861) );
and2_1 U824 ( .Z(N3688), .A(N210), .B(N2861) );
and2_1 U825 ( .Z(N3689), .A(N206), .B(N2861) );
inv_1 U826 ( .Z(N3691), .A(N2891) );
or2_1 U827 ( .Z(N3700), .A(N2907), .B(N3444) );
or2_1 U828 ( .Z(N3701), .A(N2908), .B(N3445) );
or2_1 U829 ( .Z(N3702), .A(N2909), .B(N3446) );
or3_1 U830 ( .Z(N3703), .A(N2911), .B(N3448), .C(N479) );
or3_1 U831 ( .Z(N3704), .A(N2912), .B(N3449), .C(N490) );
or2_1 U832 ( .Z(N3705), .A(N2910), .B(N3447) );
or2_1 U833 ( .Z(N3708), .A(N2919), .B(N3450) );
or2_1 U834 ( .Z(N3709), .A(N2921), .B(N3451) );
or2_1 U835 ( .Z(N3710), .A(N2922), .B(N3452) );
or3_1 U836 ( .Z(N3711), .A(N2923), .B(N3453), .C(N503) );
or3_1 U837 ( .Z(N3712), .A(N2924), .B(N3454), .C(N523) );
or3_1 U838 ( .Z(N3713), .A(N2925), .B(N3455), .C(N534) );
or2_1 U839 ( .Z(N3715), .A(N2934), .B(N3459) );
or2_1 U840 ( .Z(N3716), .A(N2935), .B(N3460) );
or2_1 U841 ( .Z(N3717), .A(N2936), .B(N3461) );
or2_1 U842 ( .Z(N3718), .A(N2937), .B(N3462) );
or3_1 U843 ( .Z(N3719), .A(N2938), .B(N3463), .C(N389) );
or3_1 U844 ( .Z(N3720), .A(N2939), .B(N3464), .C(N400) );
or3_1 U845 ( .Z(N3721), .A(N2940), .B(N3465), .C(N411) );
or3_1 U846 ( .Z(N3722), .A(N2941), .B(N3466), .C(N374) );
and2_1 U847 ( .Z(N3723), .A(N369), .B(N2942) );
and2_1 U848 ( .Z(N3724), .A(N361), .B(N2942) );
and2_1 U849 ( .Z(N3725), .A(N351), .B(N2942) );
and2_1 U850 ( .Z(N3726), .A(N341), .B(N2942) );
and2_1 U851 ( .Z(N3727), .A(N324), .B(N2948) );
and2_1 U852 ( .Z(N3728), .A(N316), .B(N2948) );
and2_1 U853 ( .Z(N3729), .A(N308), .B(N2948) );
and2_1 U854 ( .Z(N3730), .A(N302), .B(N2948) );
and2_1 U855 ( .Z(N3731), .A(N293), .B(N2948) );
or2_1 U856 ( .Z(N3732), .A(N2942), .B(N2958) );
and2_1 U857 ( .Z(N3738), .A(N83), .B(N2964) );
and2_1 U858 ( .Z(N3739), .A(N87), .B(N2964) );
and2_1 U859 ( .Z(N3740), .A(N34), .B(N2964) );
and2_1 U860 ( .Z(N3741), .A(N34), .B(N2964) );
or2_1 U861 ( .Z(N3742), .A(N2979), .B(N3481) );
or2_1 U862 ( .Z(N3743), .A(N2981), .B(N3483) );
or2_1 U863 ( .Z(N3744), .A(N2982), .B(N3484) );
or3_1 U864 ( .Z(N3745), .A(N2983), .B(N3485), .C(N503) );
or3_1 U865 ( .Z(N3746), .A(N2985), .B(N3486), .C(N523) );
or3_1 U866 ( .Z(N3747), .A(N2986), .B(N3487), .C(N534) );
or2_1 U867 ( .Z(N3748), .A(N2993), .B(N3488) );
or2_1 U868 ( .Z(N3749), .A(N2994), .B(N3489) );
or2_1 U869 ( .Z(N3750), .A(N2995), .B(N3490) );
or3_1 U870 ( .Z(N3751), .A(N2997), .B(N3492), .C(N479) );
or3_1 U871 ( .Z(N3752), .A(N2998), .B(N3493), .C(N490) );
inv_1 U872 ( .Z(N3753), .A(N3000) );
inv_1 U873 ( .Z(N3754), .A(N3003) );
inv_1 U874 ( .Z(N3755), .A(N3007) );
inv_1 U875 ( .Z(N3756), .A(N3010) );
or2_1 U876 ( .Z(N3757), .A(N3013), .B(N3502) );
and3_1 U877 ( .Z(N3758), .A(N1315), .B(N446), .C(N3003) );
or2_1 U878 ( .Z(N3759), .A(N3014), .B(N3503) );
and3_1 U879 ( .Z(N3760), .A(N1315), .B(N446), .C(N3010) );
and2_1 U880 ( .Z(N3761), .A(N1675), .B(N3000) );
and2_1 U881 ( .Z(N3762), .A(N1675), .B(N3007) );
or2_1 U882 ( .Z(N3763), .A(N3023), .B(N3504) );
or2_1 U883 ( .Z(N3764), .A(N3024), .B(N3505) );
or2_1 U884 ( .Z(N3765), .A(N3025), .B(N3506) );
or2_1 U885 ( .Z(N3766), .A(N3026), .B(N3507) );
or3_1 U886 ( .Z(N3767), .A(N3027), .B(N3508), .C(N457) );
or3_1 U887 ( .Z(N3768), .A(N3028), .B(N3509), .C(N468) );
or3_1 U888 ( .Z(N3769), .A(N3029), .B(N3510), .C(N422) );
or3_1 U889 ( .Z(N3770), .A(N3030), .B(N3511), .C(N435) );
nand2_1 U890 ( .Z(N3771), .A(N3512), .B(N3513) );
nand2_1 U891 ( .Z(N3775), .A(N3514), .B(N3515) );
inv_1 U892 ( .Z(N3779), .A(N3035) );
inv_1 U893 ( .Z(N3780), .A(N3038) );
and3_1 U894 ( .Z(N3781), .A(N117), .B(N3097), .C(N1769) );
and3_1 U895 ( .Z(N3782), .A(N126), .B(N3097), .C(N1769) );
and3_1 U896 ( .Z(N3783), .A(N127), .B(N3097), .C(N1769) );
and3_1 U897 ( .Z(N3784), .A(N128), .B(N3097), .C(N1769) );
and3_1 U898 ( .Z(N3785), .A(N131), .B(N3119), .C(N1785) );
and3_1 U899 ( .Z(N3786), .A(N129), .B(N3119), .C(N1785) );
and3_1 U900 ( .Z(N3787), .A(N119), .B(N3119), .C(N1785) );
and3_1 U901 ( .Z(N3788), .A(N130), .B(N3119), .C(N1785) );
nand2_1 U902 ( .Z(N3789), .A(N3558), .B(N3559) );
nand2_1 U903 ( .Z(N3793), .A(N3560), .B(N3561) );
nand2_1 U904 ( .Z(N3797), .A(N3562), .B(N3563) );
and3_1 U905 ( .Z(N3800), .A(N122), .B(N3147), .C(N1800) );
and3_1 U906 ( .Z(N3801), .A(N113), .B(N3147), .C(N1800) );
and3_1 U907 ( .Z(N3802), .A(N53), .B(N3147), .C(N1800) );
and3_1 U908 ( .Z(N3803), .A(N114), .B(N3147), .C(N1800) );
and3_1 U909 ( .Z(N3804), .A(N115), .B(N3147), .C(N1800) );
and3_1 U910 ( .Z(N3805), .A(N52), .B(N3169), .C(N1814) );
and3_1 U911 ( .Z(N3806), .A(N112), .B(N3169), .C(N1814) );
and3_1 U912 ( .Z(N3807), .A(N116), .B(N3169), .C(N1814) );
and3_1 U913 ( .Z(N3808), .A(N121), .B(N3169), .C(N1814) );
and3_1 U914 ( .Z(N3809), .A(N123), .B(N3169), .C(N1814) );
nand2_1 U915 ( .Z(N3810), .A(N3607), .B(N3608) );
nand2_1 U916 ( .Z(N3813), .A(N3605), .B(N3606) );
and2_1 U917 ( .Z(N3816), .A(N3482), .B(N2984) );
or2_1 U918 ( .Z(N3819), .A(N2996), .B(N3491) );
inv_1 U919 ( .Z(N3822), .A(N3200) );
nand2_1 U920 ( .Z(N3823), .A(N3200), .B(N3203) );
nand2_1 U921 ( .Z(N3824), .A(N3609), .B(N3610) );
inv_1 U922 ( .Z(N3827), .A(N3456) );
or2_1 U923 ( .Z(N3828), .A(N3739), .B(N2970) );
or2_1 U924 ( .Z(N3829), .A(N3740), .B(N2971) );
or2_1 U925 ( .Z(N3830), .A(N3741), .B(N2972) );
or2_1 U926 ( .Z(N3831), .A(N3738), .B(N2969) );
inv_1 U927 ( .Z(N3834), .A(N3664) );
inv_1 U928 ( .Z(N3835), .A(N3665) );
inv_1 U929 ( .Z(N3836), .A(N3666) );
inv_1 U930 ( .Z(N3837), .A(N3667) );
inv_1 U931 ( .Z(N3838), .A(N3672) );
inv_1 U932 ( .Z(N3839), .A(N3673) );
inv_1 U933 ( .Z(N3840), .A(N3674) );
inv_1 U934 ( .Z(N3841), .A(N3675) );
or2_1 U935 ( .Z(N3842), .A(N3681), .B(N2868) );
or2_1 U936 ( .Z(N3849), .A(N3682), .B(N2869) );
or2_1 U937 ( .Z(N3855), .A(N3683), .B(N2870) );
or2_1 U938 ( .Z(N3861), .A(N3684), .B(N2871) );
or2_1 U939 ( .Z(N3867), .A(N3685), .B(N2872) );
or2_1 U940 ( .Z(N3873), .A(N3686), .B(N2873) );
or2_1 U941 ( .Z(N3881), .A(N3687), .B(N2874) );
or2_1 U942 ( .Z(N3887), .A(N3688), .B(N2875) );
or2_1 U943 ( .Z(N3893), .A(N3689), .B(N2876) );
inv_1 U944 ( .Z(N3908), .A(N3701) );
inv_1 U945 ( .Z(N3909), .A(N3702) );
inv_1 U946 ( .Z(N3911), .A(N3700) );
inv_1 U947 ( .Z(N3914), .A(N3708) );
inv_1 U948 ( .Z(N3915), .A(N3709) );
inv_1 U949 ( .Z(N3916), .A(N3710) );
inv_1 U950 ( .Z(N3917), .A(N3715) );
inv_1 U951 ( .Z(N3918), .A(N3716) );
inv_1 U952 ( .Z(N3919), .A(N3717) );
inv_1 U953 ( .Z(N3920), .A(N3718) );
or2_1 U954 ( .Z(N3921), .A(N3724), .B(N2955) );
or2_1 U955 ( .Z(N3927), .A(N3725), .B(N2956) );
or2_1 U956 ( .Z(N3933), .A(N3726), .B(N2957) );
or2_1 U957 ( .Z(N3942), .A(N3727), .B(N2959) );
or2_1 U958 ( .Z(N3948), .A(N3728), .B(N2960) );
or2_1 U959 ( .Z(N3956), .A(N3729), .B(N2961) );
or2_1 U960 ( .Z(N3962), .A(N3730), .B(N2962) );
or2_1 U961 ( .Z(N3968), .A(N3731), .B(N2963) );
inv_1 U962 ( .Z(N3975), .A(N3742) );
inv_1 U963 ( .Z(N3976), .A(N3743) );
inv_1 U964 ( .Z(N3977), .A(N3744) );
inv_1 U965 ( .Z(N3978), .A(N3749) );
inv_1 U966 ( .Z(N3979), .A(N3750) );
and3_1 U967 ( .Z(N3980), .A(N446), .B(N1292), .C(N3754) );
and3_1 U968 ( .Z(N3981), .A(N446), .B(N1292), .C(N3756) );
and2_1 U969 ( .Z(N3982), .A(N1271), .B(N3753) );
and2_1 U970 ( .Z(N3983), .A(N1271), .B(N3755) );
inv_1 U971 ( .Z(N3984), .A(N3757) );
inv_1 U972 ( .Z(N3987), .A(N3759) );
inv_1 U973 ( .Z(N3988), .A(N3763) );
inv_1 U974 ( .Z(N3989), .A(N3764) );
inv_1 U975 ( .Z(N3990), .A(N3765) );
inv_1 U976 ( .Z(N3991), .A(N3766) );
and3_1 U977 ( .Z(N3998), .A(N3456), .B(N3119), .C(N3130) );
or2_1 U978 ( .Z(N4008), .A(N3723), .B(N2954) );
or2_1 U979 ( .Z(N4011), .A(N3680), .B(N2867) );
inv_1 U980 ( .Z(N4021), .A(N3748) );
nand2_1 U981 ( .Z(N4024), .A(N1968), .B(N3822) );
inv_1 U982 ( .Z(N4027), .A(N3705) );
and2_1 U983 ( .Z(N4031), .A(N3828), .B(N1583) );
and3_1 U984 ( .Z(N4032), .A(N24), .B(N2882), .C(N3691) );
and3_1 U985 ( .Z(N4033), .A(N25), .B(N1482), .C(N3691) );
and3_1 U986 ( .Z(N4034), .A(N26), .B(N2882), .C(N3691) );
and3_1 U987 ( .Z(N4035), .A(N81), .B(N1482), .C(N3691) );
and2_1 U988 ( .Z(N4036), .A(N3829), .B(N1583) );
and3_1 U989 ( .Z(N4037), .A(N79), .B(N2882), .C(N3691) );
and3_1 U990 ( .Z(N4038), .A(N23), .B(N1482), .C(N3691) );
and3_1 U991 ( .Z(N4039), .A(N82), .B(N2882), .C(N3691) );
and3_1 U992 ( .Z(N4040), .A(N80), .B(N1482), .C(N3691) );
and2_1 U993 ( .Z(N4041), .A(N3830), .B(N1583) );
and2_1 U994 ( .Z(N4042), .A(N3831), .B(N1583) );
and2_1 U995 ( .Z(N4067), .A(N3732), .B(N514) );
and2_1 U996 ( .Z(N4080), .A(N514), .B(N3732) );
and2_1 U997 ( .Z(N4088), .A(N3834), .B(N3668) );
and2_1 U998 ( .Z(N4091), .A(N3835), .B(N3669) );
and2_1 U999 ( .Z(N4094), .A(N3836), .B(N3670) );
and2_1 U1000 ( .Z(N4097), .A(N3837), .B(N3671) );
and2_1 U1001 ( .Z(N4100), .A(N3838), .B(N3676) );
and2_1 U1002 ( .Z(N4103), .A(N3839), .B(N3677) );
and2_1 U1003 ( .Z(N4106), .A(N3840), .B(N3678) );
and2_1 U1004 ( .Z(N4109), .A(N3841), .B(N3679) );
and2_1 U1005 ( .Z(N4144), .A(N3908), .B(N3703) );
and2_1 U1006 ( .Z(N4147), .A(N3909), .B(N3704) );
buf_1 U1007 ( .Z(N4150), .A(N3705) );
and2_1 U1008 ( .Z(N4153), .A(N3914), .B(N3711) );
and2_1 U1009 ( .Z(N4156), .A(N3915), .B(N3712) );
and2_1 U1010 ( .Z(N4159), .A(N3916), .B(N3713) );
or2_1 U1011 ( .Z(N4183), .A(N3758), .B(N3980) );
or2_1 U1012 ( .Z(N4184), .A(N3760), .B(N3981) );
or3_1 U1013 ( .Z(N4185), .A(N3761), .B(N3982), .C(N446) );
or3_1 U1014 ( .Z(N4186), .A(N3762), .B(N3983), .C(N446) );
inv_1 U1015 ( .Z(N4188), .A(N3771) );
inv_1 U1016 ( .Z(N4191), .A(N3775) );
and3_1 U1017 ( .Z(N4196), .A(N3775), .B(N3771), .C(N3035) );
and3_1 U1018 ( .Z(N4197), .A(N3987), .B(N3119), .C(N3130) );
and2_1 U1019 ( .Z(N4198), .A(N3920), .B(N3722) );
inv_1 U1020 ( .Z(N4199), .A(N3816) );
inv_1 U1021 ( .Z(N4200), .A(N3789) );
inv_1 U1022 ( .Z(N4203), .A(N3793) );
buf_1 U1023 ( .Z(N4206), .A(N3797) );
buf_1 U1024 ( .Z(N4209), .A(N3797) );
buf_1 U1025 ( .Z(N4212), .A(N3732) );
buf_1 U1026 ( .Z(N4215), .A(N3732) );
buf_1 U1027 ( .Z(N4219), .A(N3732) );
inv_1 U1028 ( .Z(N4223), .A(N3810) );
inv_1 U1029 ( .Z(N4224), .A(N3813) );
and2_1 U1030 ( .Z(N4225), .A(N3918), .B(N3720) );
and2_1 U1031 ( .Z(N4228), .A(N3919), .B(N3721) );
and2_1 U1032 ( .Z(N4231), .A(N3991), .B(N3770) );
and2_1 U1033 ( .Z(N4234), .A(N3917), .B(N3719) );
and2_1 U1034 ( .Z(N4237), .A(N3989), .B(N3768) );
and2_1 U1035 ( .Z(N4240), .A(N3990), .B(N3769) );
and2_1 U1036 ( .Z(N4243), .A(N3988), .B(N3767) );
and2_1 U1037 ( .Z(N4246), .A(N3976), .B(N3746) );
and2_1 U1038 ( .Z(N4249), .A(N3977), .B(N3747) );
and2_1 U1039 ( .Z(N4252), .A(N3975), .B(N3745) );
and2_1 U1040 ( .Z(N4255), .A(N3978), .B(N3751) );
and2_1 U1041 ( .Z(N4258), .A(N3979), .B(N3752) );
inv_1 U1042 ( .Z(N4263), .A(N3819) );
nand2_1 U1043 ( .Z(N4264), .A(N4024), .B(N3823) );
inv_1 U1044 ( .Z(N4267), .A(N3824) );
and2_1 U1045 ( .Z(N4268), .A(N446), .B(N3893) );
inv_1 U1046 ( .Z(N4269), .A(N3911) );
inv_1 U1047 ( .Z(N4270), .A(N3984) );
and2_1 U1048 ( .Z(N4271), .A(N3893), .B(N446) );
inv_1 U1049 ( .Z(N4272), .A(N4031) );
or4_1 U1050 ( .Z(N4273), .A(N4032), .B(N4033), .C(N3614), .D(N3615) );
or4_1 U1051 ( .Z(N4274), .A(N4034), .B(N4035), .C(N3625), .D(N3626) );
inv_1 U1052 ( .Z(N4275), .A(N4036) );
or4_1 U1053 ( .Z(N4276), .A(N4037), .B(N4038), .C(N3636), .D(N3637) );
or4_1 U1054 ( .Z(N4277), .A(N4039), .B(N4040), .C(N3639), .D(N3640) );
inv_1 U1055 ( .Z(N4278), .A(N4041) );
inv_1 U1056 ( .Z(N4279), .A(N4042) );
and2_1 U1057 ( .Z(N4280), .A(N3887), .B(N457) );
and2_1 U1058 ( .Z(N4284), .A(N3881), .B(N468) );
and2_1 U1059 ( .Z(N4290), .A(N422), .B(N3873) );
and2_1 U1060 ( .Z(N4297), .A(N3867), .B(N435) );
and2_1 U1061 ( .Z(N4298), .A(N3861), .B(N389) );
and2_1 U1062 ( .Z(N4301), .A(N3855), .B(N400) );
and2_1 U1063 ( .Z(N4305), .A(N3849), .B(N411) );
and2_1 U1064 ( .Z(N4310), .A(N3842), .B(N374) );
and2_1 U1065 ( .Z(N4316), .A(N457), .B(N3887) );
and2_1 U1066 ( .Z(N4320), .A(N468), .B(N3881) );
and2_1 U1067 ( .Z(N4325), .A(N422), .B(N3873) );
and2_1 U1068 ( .Z(N4331), .A(N435), .B(N3867) );
and2_1 U1069 ( .Z(N4332), .A(N389), .B(N3861) );
and2_1 U1070 ( .Z(N4336), .A(N400), .B(N3855) );
and2_1 U1071 ( .Z(N4342), .A(N411), .B(N3849) );
and2_1 U1072 ( .Z(N4349), .A(N374), .B(N3842) );
inv_1 U1073 ( .Z(N4357), .A(N3968) );
inv_1 U1074 ( .Z(N4364), .A(N3962) );
buf_1 U1075 ( .Z(N4375), .A(N3962) );
and2_1 U1076 ( .Z(N4379), .A(N3956), .B(N479) );
and2_1 U1077 ( .Z(N4385), .A(N490), .B(N3948) );
and2_1 U1078 ( .Z(N4392), .A(N3942), .B(N503) );
and2_1 U1079 ( .Z(N4396), .A(N3933), .B(N523) );
and2_1 U1080 ( .Z(N4400), .A(N3927), .B(N534) );
inv_1 U1081 ( .Z(N4405), .A(N3921) );
buf_1 U1082 ( .Z(N4412), .A(N3921) );
inv_1 U1083 ( .Z(N4418), .A(N3968) );
inv_1 U1084 ( .Z(N4425), .A(N3962) );
buf_1 U1085 ( .Z(N4436), .A(N3962) );
and2_1 U1086 ( .Z(N4440), .A(N479), .B(N3956) );
and2_1 U1087 ( .Z(N4445), .A(N490), .B(N3948) );
and2_1 U1088 ( .Z(N4451), .A(N503), .B(N3942) );
and2_1 U1089 ( .Z(N4456), .A(N523), .B(N3933) );
and2_1 U1090 ( .Z(N4462), .A(N534), .B(N3927) );
buf_1 U1091 ( .Z(N4469), .A(N3921) );
inv_1 U1092 ( .Z(N4477), .A(N3921) );
buf_1 U1093 ( .Z(N4512), .A(N3968) );
inv_1 U1094 ( .Z(N4515), .A(N4183) );
inv_1 U1095 ( .Z(N4516), .A(N4184) );
inv_1 U1096 ( .Z(N4521), .A(N4008) );
inv_1 U1097 ( .Z(N4523), .A(N4011) );
inv_1 U1098 ( .Z(N4524), .A(N4198) );
inv_1 U1099 ( .Z(N4532), .A(N3984) );
and3_1 U1100 ( .Z(N4547), .A(N3911), .B(N3169), .C(N3180) );
buf_1 U1101 ( .Z(N4548), .A(N3893) );
buf_1 U1102 ( .Z(N4551), .A(N3887) );
buf_1 U1103 ( .Z(N4554), .A(N3881) );
buf_1 U1104 ( .Z(N4557), .A(N3873) );
buf_1 U1105 ( .Z(N4560), .A(N3867) );
buf_1 U1106 ( .Z(N4563), .A(N3861) );
buf_1 U1107 ( .Z(N4566), .A(N3855) );
buf_1 U1108 ( .Z(N4569), .A(N3849) );
buf_1 U1109 ( .Z(N4572), .A(N3842) );
nor2_1 U1110 ( .Z(N4575), .A(N422), .B(N3873) );
buf_1 U1111 ( .Z(N4578), .A(N3893) );
buf_1 U1112 ( .Z(N4581), .A(N3887) );
buf_1 U1113 ( .Z(N4584), .A(N3881) );
buf_1 U1114 ( .Z(N4587), .A(N3867) );
buf_1 U1115 ( .Z(N4590), .A(N3861) );
buf_1 U1116 ( .Z(N4593), .A(N3855) );
buf_1 U1117 ( .Z(N4596), .A(N3849) );
buf_1 U1118 ( .Z(N4599), .A(N3873) );
buf_1 U1119 ( .Z(N4602), .A(N3842) );
nor2_1 U1120 ( .Z(N4605), .A(N422), .B(N3873) );
nor2_1 U1121 ( .Z(N4608), .A(N374), .B(N3842) );
buf_1 U1122 ( .Z(N4611), .A(N3956) );
buf_1 U1123 ( .Z(N4614), .A(N3948) );
buf_1 U1124 ( .Z(N4617), .A(N3942) );
buf_1 U1125 ( .Z(N4621), .A(N3933) );
buf_1 U1126 ( .Z(N4624), .A(N3927) );
nor2_1 U1127 ( .Z(N4627), .A(N490), .B(N3948) );
buf_1 U1128 ( .Z(N4630), .A(N3956) );
buf_1 U1129 ( .Z(N4633), .A(N3942) );
buf_1 U1130 ( .Z(N4637), .A(N3933) );
buf_1 U1131 ( .Z(N4640), .A(N3927) );
buf_1 U1132 ( .Z(N4643), .A(N3948) );
nor2_1 U1133 ( .Z(N4646), .A(N490), .B(N3948) );
buf_1 U1134 ( .Z(N4649), .A(N3927) );
buf_1 U1135 ( .Z(N4652), .A(N3933) );
buf_1 U1136 ( .Z(N4655), .A(N3921) );
buf_1 U1137 ( .Z(N4658), .A(N3942) );
buf_1 U1138 ( .Z(N4662), .A(N3956) );
buf_1 U1139 ( .Z(N4665), .A(N3948) );
buf_1 U1140 ( .Z(N4668), .A(N3968) );
buf_1 U1141 ( .Z(N4671), .A(N3962) );
buf_1 U1142 ( .Z(N4674), .A(N3873) );
buf_1 U1143 ( .Z(N4677), .A(N3867) );
buf_1 U1144 ( .Z(N4680), .A(N3887) );
buf_1 U1145 ( .Z(N4683), .A(N3881) );
buf_1 U1146 ( .Z(N4686), .A(N3893) );
buf_1 U1147 ( .Z(N4689), .A(N3849) );
buf_1 U1148 ( .Z(N4692), .A(N3842) );
buf_1 U1149 ( .Z(N4695), .A(N3861) );
buf_1 U1150 ( .Z(N4698), .A(N3855) );
nand2_1 U1151 ( .Z(N4701), .A(N3813), .B(N4223) );
nand2_1 U1152 ( .Z(N4702), .A(N3810), .B(N4224) );
inv_1 U1153 ( .Z(N4720), .A(N4021) );
nand2_1 U1154 ( .Z(N4721), .A(N4021), .B(N4263) );
inv_1 U1155 ( .Z(N4724), .A(N4147) );
inv_1 U1156 ( .Z(N4725), .A(N4144) );
inv_1 U1157 ( .Z(N4726), .A(N4159) );
inv_1 U1158 ( .Z(N4727), .A(N4156) );
inv_1 U1159 ( .Z(N4728), .A(N4153) );
inv_1 U1160 ( .Z(N4729), .A(N4097) );
inv_1 U1161 ( .Z(N4730), .A(N4094) );
inv_1 U1162 ( .Z(N4731), .A(N4091) );
inv_1 U1163 ( .Z(N4732), .A(N4088) );
inv_1 U1164 ( .Z(N4733), .A(N4109) );
inv_1 U1165 ( .Z(N4734), .A(N4106) );
inv_1 U1166 ( .Z(N4735), .A(N4103) );
inv_1 U1167 ( .Z(N4736), .A(N4100) );
and2_1 U1168 ( .Z(N4737), .A(N4273), .B(N2877) );
and2_1 U1169 ( .Z(N4738), .A(N4274), .B(N2877) );
and2_1 U1170 ( .Z(N4739), .A(N4276), .B(N2877) );
and2_1 U1171 ( .Z(N4740), .A(N4277), .B(N2877) );
and3_1 U1172 ( .Z(N4741), .A(N4150), .B(N1758), .C(N1755) );
inv_1 U1173 ( .Z(N4855), .A(N4212) );
nand2_1 U1174 ( .Z(N4856), .A(N4212), .B(N2712) );
nand2_1 U1175 ( .Z(N4908), .A(N4215), .B(N2718) );
inv_1 U1176 ( .Z(N4909), .A(N4215) );
and2_1 U1177 ( .Z(N4939), .A(N4515), .B(N4185) );
and2_1 U1178 ( .Z(N4942), .A(N4516), .B(N4186) );
inv_1 U1179 ( .Z(N4947), .A(N4219) );
and3_1 U1180 ( .Z(N4953), .A(N4188), .B(N3775), .C(N3779) );
and3_1 U1181 ( .Z(N4954), .A(N3771), .B(N4191), .C(N3780) );
and3_1 U1182 ( .Z(N4955), .A(N4191), .B(N4188), .C(N3038) );
and3_1 U1183 ( .Z(N4956), .A(N4109), .B(N3097), .C(N3108) );
and3_1 U1184 ( .Z(N4957), .A(N4106), .B(N3097), .C(N3108) );
and3_1 U1185 ( .Z(N4958), .A(N4103), .B(N3097), .C(N3108) );
and3_1 U1186 ( .Z(N4959), .A(N4100), .B(N3097), .C(N3108) );
and3_1 U1187 ( .Z(N4960), .A(N4159), .B(N3119), .C(N3130) );
and3_1 U1188 ( .Z(N4961), .A(N4156), .B(N3119), .C(N3130) );
inv_1 U1189 ( .Z(N4965), .A(N4225) );
inv_1 U1190 ( .Z(N4966), .A(N4228) );
inv_1 U1191 ( .Z(N4967), .A(N4231) );
inv_1 U1192 ( .Z(N4968), .A(N4234) );
inv_1 U1193 ( .Z(N4972), .A(N4246) );
inv_1 U1194 ( .Z(N4973), .A(N4249) );
inv_1 U1195 ( .Z(N4974), .A(N4252) );
nand2_1 U1196 ( .Z(N4975), .A(N4252), .B(N4199) );
inv_1 U1197 ( .Z(N4976), .A(N4206) );
inv_1 U1198 ( .Z(N4977), .A(N4209) );
and3_1 U1199 ( .Z(N4978), .A(N3793), .B(N3789), .C(N4206) );
and3_1 U1200 ( .Z(N4979), .A(N4203), .B(N4200), .C(N4209) );
and3_1 U1201 ( .Z(N4980), .A(N4097), .B(N3147), .C(N3158) );
and3_1 U1202 ( .Z(N4981), .A(N4094), .B(N3147), .C(N3158) );
and3_1 U1203 ( .Z(N4982), .A(N4091), .B(N3147), .C(N3158) );
and3_1 U1204 ( .Z(N4983), .A(N4088), .B(N3147), .C(N3158) );
and3_1 U1205 ( .Z(N4984), .A(N4153), .B(N3169), .C(N3180) );
and3_1 U1206 ( .Z(N4985), .A(N4147), .B(N3169), .C(N3180) );
and3_1 U1207 ( .Z(N4986), .A(N4144), .B(N3169), .C(N3180) );
and3_1 U1208 ( .Z(N4987), .A(N4150), .B(N3169), .C(N3180) );
nand2_1 U1209 ( .Z(N5049), .A(N4701), .B(N4702) );
inv_1 U1210 ( .Z(N5052), .A(N4237) );
inv_1 U1211 ( .Z(N5053), .A(N4240) );
inv_1 U1212 ( .Z(N5054), .A(N4243) );
inv_1 U1213 ( .Z(N5055), .A(N4255) );
inv_1 U1214 ( .Z(N5056), .A(N4258) );
nand2_1 U1215 ( .Z(N5057), .A(N3819), .B(N4720) );
inv_1 U1216 ( .Z(N5058), .A(N4264) );
nand2_1 U1217 ( .Z(N5059), .A(N4264), .B(N4267) );
and4_1 U1218 ( .Z(N5060), .A(N4724), .B(N4725), .C(N4269), .D(N4027) );
and4_1 U1219 ( .Z(N5061), .A(N4726), .B(N4727), .C(N3827), .D(N4728) );
and4_1 U1220 ( .Z(N5062), .A(N4729), .B(N4730), .C(N4731), .D(N4732) );
and4_1 U1221 ( .Z(N5063), .A(N4733), .B(N4734), .C(N4735), .D(N4736) );
and2_1 U1222 ( .Z(N5065), .A(N4357), .B(N4375) );
and3_1 U1223 ( .Z(N5066), .A(N4364), .B(N4357), .C(N4379) );
and2_1 U1224 ( .Z(N5067), .A(N4418), .B(N4436) );
and3_1 U1225 ( .Z(N5068), .A(N4425), .B(N4418), .C(N4440) );
inv_1 U1226 ( .Z(N5069), .A(N4548) );
nand2_1 U1227 ( .Z(N5070), .A(N4548), .B(N2628) );
inv_1 U1228 ( .Z(N5071), .A(N4551) );
nand2_1 U1229 ( .Z(N5072), .A(N4551), .B(N2629) );
inv_1 U1230 ( .Z(N5073), .A(N4554) );
nand2_1 U1231 ( .Z(N5074), .A(N4554), .B(N2630) );
inv_1 U1232 ( .Z(N5075), .A(N4557) );
nand2_1 U1233 ( .Z(N5076), .A(N4557), .B(N2631) );
inv_1 U1234 ( .Z(N5077), .A(N4560) );
nand2_1 U1235 ( .Z(N5078), .A(N4560), .B(N2632) );
inv_1 U1236 ( .Z(N5079), .A(N4563) );
nand2_1 U1237 ( .Z(N5080), .A(N4563), .B(N2633) );
inv_1 U1238 ( .Z(N5081), .A(N4566) );
nand2_1 U1239 ( .Z(N5082), .A(N4566), .B(N2634) );
inv_1 U1240 ( .Z(N5083), .A(N4569) );
nand2_1 U1241 ( .Z(N5084), .A(N4569), .B(N2635) );
inv_1 U1242 ( .Z(N5085), .A(N4572) );
nand2_1 U1243 ( .Z(N5086), .A(N4572), .B(N2636) );
inv_1 U1244 ( .Z(N5087), .A(N4575) );
nand2_1 U1245 ( .Z(N5088), .A(N4578), .B(N2638) );
inv_1 U1246 ( .Z(N5089), .A(N4578) );
nand2_1 U1247 ( .Z(N5090), .A(N4581), .B(N2639) );
inv_1 U1248 ( .Z(N5091), .A(N4581) );
nand2_1 U1249 ( .Z(N5092), .A(N4584), .B(N2640) );
inv_1 U1250 ( .Z(N5093), .A(N4584) );
nand2_1 U1251 ( .Z(N5094), .A(N4587), .B(N2641) );
inv_1 U1252 ( .Z(N5095), .A(N4587) );
nand2_1 U1253 ( .Z(N5096), .A(N4590), .B(N2642) );
inv_1 U1254 ( .Z(N5097), .A(N4590) );
nand2_1 U1255 ( .Z(N5098), .A(N4593), .B(N2643) );
inv_1 U1256 ( .Z(N5099), .A(N4593) );
nand2_1 U1257 ( .Z(N5100), .A(N4596), .B(N2644) );
inv_1 U1258 ( .Z(N5101), .A(N4596) );
nand2_1 U1259 ( .Z(N5102), .A(N4599), .B(N2645) );
inv_1 U1260 ( .Z(N5103), .A(N4599) );
nand2_1 U1261 ( .Z(N5104), .A(N4602), .B(N2646) );
inv_1 U1262 ( .Z(N5105), .A(N4602) );
inv_1 U1263 ( .Z(N5106), .A(N4611) );
nand2_1 U1264 ( .Z(N5107), .A(N4611), .B(N2709) );
inv_1 U1265 ( .Z(N5108), .A(N4614) );
nand2_1 U1266 ( .Z(N5109), .A(N4614), .B(N2710) );
inv_1 U1267 ( .Z(N5110), .A(N4617) );
nand2_1 U1268 ( .Z(N5111), .A(N4617), .B(N2711) );
nand2_1 U1269 ( .Z(N5112), .A(N1890), .B(N4855) );
inv_1 U1270 ( .Z(N5113), .A(N4621) );
nand2_1 U1271 ( .Z(N5114), .A(N4621), .B(N2713) );
inv_1 U1272 ( .Z(N5115), .A(N4624) );
nand2_1 U1273 ( .Z(N5116), .A(N4624), .B(N2714) );
and2_1 U1274 ( .Z(N5117), .A(N4364), .B(N4379) );
and2_1 U1275 ( .Z(N5118), .A(N4364), .B(N4379) );
and2_1 U1276 ( .Z(N5119), .A(N54), .B(N4405) );
inv_1 U1277 ( .Z(N5120), .A(N4627) );
nand2_1 U1278 ( .Z(N5121), .A(N4630), .B(N2716) );
inv_1 U1279 ( .Z(N5122), .A(N4630) );
nand2_1 U1280 ( .Z(N5123), .A(N4633), .B(N2717) );
inv_1 U1281 ( .Z(N5124), .A(N4633) );
nand2_1 U1282 ( .Z(N5125), .A(N1908), .B(N4909) );
nand2_1 U1283 ( .Z(N5126), .A(N4637), .B(N2719) );
inv_1 U1284 ( .Z(N5127), .A(N4637) );
nand2_1 U1285 ( .Z(N5128), .A(N4640), .B(N2720) );
inv_1 U1286 ( .Z(N5129), .A(N4640) );
nand2_1 U1287 ( .Z(N5130), .A(N4643), .B(N2721) );
inv_1 U1288 ( .Z(N5131), .A(N4643) );
and2_1 U1289 ( .Z(N5132), .A(N4425), .B(N4440) );
and2_1 U1290 ( .Z(N5133), .A(N4425), .B(N4440) );
inv_1 U1291 ( .Z(N5135), .A(N4649) );
inv_1 U1292 ( .Z(N5136), .A(N4652) );
nand2_1 U1293 ( .Z(N5137), .A(N4655), .B(N4521) );
inv_1 U1294 ( .Z(N5138), .A(N4655) );
inv_1 U1295 ( .Z(N5139), .A(N4658) );
nand2_1 U1296 ( .Z(N5140), .A(N4658), .B(N4947) );
inv_1 U1297 ( .Z(N5141), .A(N4674) );
inv_1 U1298 ( .Z(N5142), .A(N4677) );
inv_1 U1299 ( .Z(N5143), .A(N4680) );
inv_1 U1300 ( .Z(N5144), .A(N4683) );
nand2_1 U1301 ( .Z(N5145), .A(N4686), .B(N4523) );
inv_1 U1302 ( .Z(N5146), .A(N4686) );
nor2_1 U1303 ( .Z(N5147), .A(N4953), .B(N4196) );
nor2_1 U1304 ( .Z(N5148), .A(N4954), .B(N4955) );
inv_1 U1305 ( .Z(N5150), .A(N4524) );
nand2_1 U1306 ( .Z(N5153), .A(N4228), .B(N4965) );
nand2_1 U1307 ( .Z(N5154), .A(N4225), .B(N4966) );
nand2_1 U1308 ( .Z(N5155), .A(N4234), .B(N4967) );
nand2_1 U1309 ( .Z(N5156), .A(N4231), .B(N4968) );
inv_1 U1310 ( .Z(N5157), .A(N4532) );
nand2_1 U1311 ( .Z(N5160), .A(N4249), .B(N4972) );
nand2_1 U1312 ( .Z(N5161), .A(N4246), .B(N4973) );
nand2_1 U1313 ( .Z(N5162), .A(N3816), .B(N4974) );
and3_1 U1314 ( .Z(N5163), .A(N4200), .B(N3793), .C(N4976) );
and3_1 U1315 ( .Z(N5164), .A(N3789), .B(N4203), .C(N4977) );
and3_1 U1316 ( .Z(N5165), .A(N4942), .B(N3147), .C(N3158) );
inv_1 U1317 ( .Z(N5166), .A(N4512) );
buf_1 U1318 ( .Z(N5169), .A(N4290) );
inv_1 U1319 ( .Z(N5172), .A(N4605) );
buf_1 U1320 ( .Z(N5173), .A(N4325) );
inv_1 U1321 ( .Z(N5176), .A(N4608) );
buf_1 U1322 ( .Z(N5177), .A(N4349) );
buf_1 U1323 ( .Z(N5180), .A(N4405) );
buf_1 U1324 ( .Z(N5183), .A(N4357) );
buf_1 U1325 ( .Z(N5186), .A(N4357) );
buf_1 U1326 ( .Z(N5189), .A(N4364) );
buf_1 U1327 ( .Z(N5192), .A(N4364) );
buf_1 U1328 ( .Z(N5195), .A(N4385) );
inv_1 U1329 ( .Z(N5198), .A(N4646) );
buf_1 U1330 ( .Z(N5199), .A(N4418) );
buf_1 U1331 ( .Z(N5202), .A(N4425) );
buf_1 U1332 ( .Z(N5205), .A(N4445) );
buf_1 U1333 ( .Z(N5208), .A(N4418) );
buf_1 U1334 ( .Z(N5211), .A(N4425) );
buf_1 U1335 ( .Z(N5214), .A(N4477) );
buf_1 U1336 ( .Z(N5217), .A(N4469) );
buf_1 U1337 ( .Z(N5220), .A(N4477) );
inv_1 U1338 ( .Z(N5223), .A(N4662) );
inv_1 U1339 ( .Z(N5224), .A(N4665) );
inv_1 U1340 ( .Z(N5225), .A(N4668) );
inv_1 U1341 ( .Z(N5226), .A(N4671) );
inv_1 U1342 ( .Z(N5227), .A(N4689) );
inv_1 U1343 ( .Z(N5228), .A(N4692) );
inv_1 U1344 ( .Z(N5229), .A(N4695) );
inv_1 U1345 ( .Z(N5230), .A(N4698) );
nand2_1 U1346 ( .Z(N5232), .A(N4240), .B(N5052) );
nand2_1 U1347 ( .Z(N5233), .A(N4237), .B(N5053) );
nand2_1 U1348 ( .Z(N5234), .A(N4258), .B(N5055) );
nand2_1 U1349 ( .Z(N5235), .A(N4255), .B(N5056) );
nand2_1 U1350 ( .Z(N5236), .A(N4721), .B(N5057) );
nand2_1 U1351 ( .Z(N5239), .A(N3824), .B(N5058) );
and3_1 U1352 ( .Z(N5240), .A(N5060), .B(N5061), .C(N4270) );
inv_1 U1353 ( .Z(N5241), .A(N4939) );
nand2_1 U1354 ( .Z(N5242), .A(N1824), .B(N5069) );
nand2_1 U1355 ( .Z(N5243), .A(N1827), .B(N5071) );
nand2_1 U1356 ( .Z(N5244), .A(N1830), .B(N5073) );
nand2_1 U1357 ( .Z(N5245), .A(N1833), .B(N5075) );
nand2_1 U1358 ( .Z(N5246), .A(N1836), .B(N5077) );
nand2_1 U1359 ( .Z(N5247), .A(N1839), .B(N5079) );
nand2_1 U1360 ( .Z(N5248), .A(N1842), .B(N5081) );
nand2_1 U1361 ( .Z(N5249), .A(N1845), .B(N5083) );
nand2_1 U1362 ( .Z(N5250), .A(N1848), .B(N5085) );
nand2_1 U1363 ( .Z(N5252), .A(N1854), .B(N5089) );
nand2_1 U1364 ( .Z(N5253), .A(N1857), .B(N5091) );
nand2_1 U1365 ( .Z(N5254), .A(N1860), .B(N5093) );
nand2_1 U1366 ( .Z(N5255), .A(N1863), .B(N5095) );
nand2_1 U1367 ( .Z(N5256), .A(N1866), .B(N5097) );
nand2_1 U1368 ( .Z(N5257), .A(N1869), .B(N5099) );
nand2_1 U1369 ( .Z(N5258), .A(N1872), .B(N5101) );
nand2_1 U1370 ( .Z(N5259), .A(N1875), .B(N5103) );
nand2_1 U1371 ( .Z(N5260), .A(N1878), .B(N5105) );
nand2_1 U1372 ( .Z(N5261), .A(N1881), .B(N5106) );
nand2_1 U1373 ( .Z(N5262), .A(N1884), .B(N5108) );
nand2_1 U1374 ( .Z(N5263), .A(N1887), .B(N5110) );
nand2_1 U1375 ( .Z(N5264), .A(N5112), .B(N4856) );
nand2_1 U1376 ( .Z(N5274), .A(N1893), .B(N5113) );
nand2_1 U1377 ( .Z(N5275), .A(N1896), .B(N5115) );
nand2_1 U1378 ( .Z(N5282), .A(N1902), .B(N5122) );
nand2_1 U1379 ( .Z(N5283), .A(N1905), .B(N5124) );
nand2_1 U1380 ( .Z(N5284), .A(N4908), .B(N5125) );
nand2_1 U1381 ( .Z(N5298), .A(N1911), .B(N5127) );
nand2_1 U1382 ( .Z(N5299), .A(N1914), .B(N5129) );
nand2_1 U1383 ( .Z(N5300), .A(N1917), .B(N5131) );
nand2_1 U1384 ( .Z(N5303), .A(N4652), .B(N5135) );
nand2_1 U1385 ( .Z(N5304), .A(N4649), .B(N5136) );
nand2_1 U1386 ( .Z(N5305), .A(N4008), .B(N5138) );
nand2_1 U1387 ( .Z(N5306), .A(N4219), .B(N5139) );
nand2_1 U1388 ( .Z(N5307), .A(N4677), .B(N5141) );
nand2_1 U1389 ( .Z(N5308), .A(N4674), .B(N5142) );
nand2_1 U1390 ( .Z(N5309), .A(N4683), .B(N5143) );
nand2_1 U1391 ( .Z(N5310), .A(N4680), .B(N5144) );
nand2_1 U1392 ( .Z(N5311), .A(N4011), .B(N5146) );
inv_1 U1393 ( .Z(N5312), .A(N5049) );
nand2_1 U1394 ( .Z(N5315), .A(N5153), .B(N5154) );
nand2_1 U1395 ( .Z(N5319), .A(N5155), .B(N5156) );
nand2_1 U1396 ( .Z(N5324), .A(N5160), .B(N5161) );
nand2_1 U1397 ( .Z(N5328), .A(N5162), .B(N4975) );
nor2_1 U1398 ( .Z(N5331), .A(N5163), .B(N4978) );
nor2_1 U1399 ( .Z(N5332), .A(N5164), .B(N4979) );
or2_1 U1400 ( .Z(N5346), .A(N4412), .B(N5119) );
nand2_1 U1401 ( .Z(N5363), .A(N4665), .B(N5223) );
nand2_1 U1402 ( .Z(N5364), .A(N4662), .B(N5224) );
nand2_1 U1403 ( .Z(N5365), .A(N4671), .B(N5225) );
nand2_1 U1404 ( .Z(N5366), .A(N4668), .B(N5226) );
nand2_1 U1405 ( .Z(N5367), .A(N4692), .B(N5227) );
nand2_1 U1406 ( .Z(N5368), .A(N4689), .B(N5228) );
nand2_1 U1407 ( .Z(N5369), .A(N4698), .B(N5229) );
nand2_1 U1408 ( .Z(N5370), .A(N4695), .B(N5230) );
nand2_1 U1409 ( .Z(N5371), .A(N5148), .B(N5147) );
buf_1 U1410 ( .Z(N5374), .A(N4939) );
nand2_1 U1411 ( .Z(N5377), .A(N5232), .B(N5233) );
nand2_1 U1412 ( .Z(N5382), .A(N5234), .B(N5235) );
nand2_1 U1413 ( .Z(N5385), .A(N5239), .B(N5059) );
and3_1 U1414 ( .Z(N5388), .A(N5062), .B(N5063), .C(N5241) );
nand2_1 U1415 ( .Z(N5389), .A(N5242), .B(N5070) );
nand2_1 U1416 ( .Z(N5396), .A(N5243), .B(N5072) );
nand2_1 U1417 ( .Z(N5407), .A(N5244), .B(N5074) );
nand2_1 U1418 ( .Z(N5418), .A(N5245), .B(N5076) );
nand2_1 U1419 ( .Z(N5424), .A(N5246), .B(N5078) );
nand2_1 U1420 ( .Z(N5431), .A(N5247), .B(N5080) );
nand2_1 U1421 ( .Z(N5441), .A(N5248), .B(N5082) );
nand2_1 U1422 ( .Z(N5452), .A(N5249), .B(N5084) );
nand2_1 U1423 ( .Z(N5462), .A(N5250), .B(N5086) );
inv_1 U1424 ( .Z(N5469), .A(N5169) );
nand2_1 U1425 ( .Z(N5470), .A(N5088), .B(N5252) );
nand2_1 U1426 ( .Z(N5477), .A(N5090), .B(N5253) );
nand2_1 U1427 ( .Z(N5488), .A(N5092), .B(N5254) );
nand2_1 U1428 ( .Z(N5498), .A(N5094), .B(N5255) );
nand2_1 U1429 ( .Z(N5506), .A(N5096), .B(N5256) );
nand2_1 U1430 ( .Z(N5520), .A(N5098), .B(N5257) );
nand2_1 U1431 ( .Z(N5536), .A(N5100), .B(N5258) );
nand2_1 U1432 ( .Z(N5549), .A(N5102), .B(N5259) );
nand2_1 U1433 ( .Z(N5555), .A(N5104), .B(N5260) );
nand2_1 U1434 ( .Z(N5562), .A(N5261), .B(N5107) );
nand2_1 U1435 ( .Z(N5573), .A(N5262), .B(N5109) );
nand2_1 U1436 ( .Z(N5579), .A(N5263), .B(N5111) );
nand2_1 U1437 ( .Z(N5595), .A(N5274), .B(N5114) );
nand2_1 U1438 ( .Z(N5606), .A(N5275), .B(N5116) );
nand2_1 U1439 ( .Z(N5616), .A(N5180), .B(N2715) );
inv_1 U1440 ( .Z(N5617), .A(N5180) );
inv_1 U1441 ( .Z(N5618), .A(N5183) );
inv_1 U1442 ( .Z(N5619), .A(N5186) );
inv_1 U1443 ( .Z(N5620), .A(N5189) );
inv_1 U1444 ( .Z(N5621), .A(N5192) );
inv_1 U1445 ( .Z(N5622), .A(N5195) );
nand2_1 U1446 ( .Z(N5624), .A(N5121), .B(N5282) );
nand2_1 U1447 ( .Z(N5634), .A(N5123), .B(N5283) );
nand2_1 U1448 ( .Z(N5655), .A(N5126), .B(N5298) );
nand2_1 U1449 ( .Z(N5671), .A(N5128), .B(N5299) );
nand2_1 U1450 ( .Z(N5684), .A(N5130), .B(N5300) );
inv_1 U1451 ( .Z(N5690), .A(N5202) );
inv_1 U1452 ( .Z(N5691), .A(N5211) );
nand2_1 U1453 ( .Z(N5692), .A(N5303), .B(N5304) );
nand2_1 U1454 ( .Z(N5696), .A(N5137), .B(N5305) );
nand2_1 U1455 ( .Z(N5700), .A(N5306), .B(N5140) );
nand2_1 U1456 ( .Z(N5703), .A(N5307), .B(N5308) );
nand2_1 U1457 ( .Z(N5707), .A(N5309), .B(N5310) );
nand2_1 U1458 ( .Z(N5711), .A(N5145), .B(N5311) );
and2_1 U1459 ( .Z(N5726), .A(N5166), .B(N4512) );
inv_1 U1460 ( .Z(N5727), .A(N5173) );
inv_1 U1461 ( .Z(N5728), .A(N5177) );
inv_1 U1462 ( .Z(N5730), .A(N5199) );
inv_1 U1463 ( .Z(N5731), .A(N5205) );
inv_1 U1464 ( .Z(N5732), .A(N5208) );
inv_1 U1465 ( .Z(N5733), .A(N5214) );
inv_1 U1466 ( .Z(N5734), .A(N5217) );
inv_1 U1467 ( .Z(N5735), .A(N5220) );
nand2_1 U1468 ( .Z(N5736), .A(N5365), .B(N5366) );
nand2_1 U1469 ( .Z(N5739), .A(N5363), .B(N5364) );
nand2_1 U1470 ( .Z(N5742), .A(N5369), .B(N5370) );
nand2_1 U1471 ( .Z(N5745), .A(N5367), .B(N5368) );
inv_1 U1472 ( .Z(N5755), .A(N5236) );
nand2_1 U1473 ( .Z(N5756), .A(N5332), .B(N5331) );
and2_1 U1474 ( .Z(N5954), .A(N5264), .B(N4396) );
nand2_1 U1475 ( .Z(N5955), .A(N1899), .B(N5617) );
inv_1 U1476 ( .Z(N5956), .A(N5346) );
and2_1 U1477 ( .Z(N6005), .A(N5284), .B(N4456) );
and2_1 U1478 ( .Z(N6006), .A(N5284), .B(N4456) );
inv_1 U1479 ( .Z(N6023), .A(N5371) );
nand2_1 U1480 ( .Z(N6024), .A(N5371), .B(N5312) );
inv_1 U1481 ( .Z(N6025), .A(N5315) );
inv_1 U1482 ( .Z(N6028), .A(N5324) );
buf_1 U1483 ( .Z(N6031), .A(N5319) );
buf_1 U1484 ( .Z(N6034), .A(N5319) );
buf_1 U1485 ( .Z(N6037), .A(N5328) );
buf_1 U1486 ( .Z(N6040), .A(N5328) );
inv_1 U1487 ( .Z(N6044), .A(N5385) );
or2_1 U1488 ( .Z(N6045), .A(N5166), .B(N5726) );
buf_1 U1489 ( .Z(N6048), .A(N5264) );
buf_1 U1490 ( .Z(N6051), .A(N5284) );
buf_1 U1491 ( .Z(N6054), .A(N5284) );
inv_1 U1492 ( .Z(N6065), .A(N5374) );
nand2_1 U1493 ( .Z(N6066), .A(N5374), .B(N5054) );
inv_1 U1494 ( .Z(N6067), .A(N5377) );
inv_1 U1495 ( .Z(N6068), .A(N5382) );
nand2_1 U1496 ( .Z(N6069), .A(N5382), .B(N5755) );
and2_1 U1497 ( .Z(N6071), .A(N5470), .B(N4316) );
and3_1 U1498 ( .Z(N6072), .A(N5477), .B(N5470), .C(N4320) );
and4_1 U1499 ( .Z(N6073), .A(N5488), .B(N5470), .C(N4325), .D(N5477) );
and4_1 U1500 ( .Z(N6074), .A(N5562), .B(N4357), .C(N4385), .D(N4364) );
and2_1 U1501 ( .Z(N6075), .A(N5389), .B(N4280) );
and3_1 U1502 ( .Z(N6076), .A(N5396), .B(N5389), .C(N4284) );
and4_1 U1503 ( .Z(N6077), .A(N5407), .B(N5389), .C(N4290), .D(N5396) );
and4_1 U1504 ( .Z(N6078), .A(N5624), .B(N4418), .C(N4445), .D(N4425) );
inv_1 U1505 ( .Z(N6079), .A(N5418) );
and4_1 U1506 ( .Z(N6080), .A(N5396), .B(N5418), .C(N5407), .D(N5389) );
and2_1 U1507 ( .Z(N6083), .A(N5396), .B(N4284) );
and3_1 U1508 ( .Z(N6084), .A(N5407), .B(N4290), .C(N5396) );
and3_1 U1509 ( .Z(N6085), .A(N5418), .B(N5407), .C(N5396) );
and2_1 U1510 ( .Z(N6086), .A(N5396), .B(N4284) );
and3_1 U1511 ( .Z(N6087), .A(N4290), .B(N5407), .C(N5396) );
and2_1 U1512 ( .Z(N6088), .A(N5407), .B(N4290) );
and2_1 U1513 ( .Z(N6089), .A(N5418), .B(N5407) );
and2_1 U1514 ( .Z(N6090), .A(N5407), .B(N4290) );
and5_1 U1515 ( .Z(N6091), .A(N5431), .B(N5462), .C(N5441), .D(N5424), .E(N5452) );
and2_1 U1516 ( .Z(N6094), .A(N5424), .B(N4298) );
and3_1 U1517 ( .Z(N6095), .A(N5431), .B(N5424), .C(N4301) );
and4_1 U1518 ( .Z(N6096), .A(N5441), .B(N5424), .C(N4305), .D(N5431) );
and5_1 U1519 ( .Z(N6097), .A(N5452), .B(N5441), .C(N5424), .D(N4310), .E(N5431) );
and2_1 U1520 ( .Z(N6098), .A(N5431), .B(N4301) );
and3_1 U1521 ( .Z(N6099), .A(N5441), .B(N4305), .C(N5431) );
and4_1 U1522 ( .Z(N6100), .A(N5452), .B(N5441), .C(N4310), .D(N5431) );
and5_1 U1523 ( .Z(N6101), .A(N4), .B(N5462), .C(N5441), .D(N5452), .E(N5431) );
and2_1 U1524 ( .Z(N6102), .A(N4305), .B(N5441) );
and3_1 U1525 ( .Z(N6103), .A(N5452), .B(N5441), .C(N4310) );
and4_1 U1526 ( .Z(N6104), .A(N4), .B(N5462), .C(N5441), .D(N5452) );
and2_1 U1527 ( .Z(N6105), .A(N5452), .B(N4310) );
and3_1 U1528 ( .Z(N6106), .A(N4), .B(N5462), .C(N5452) );
and2_1 U1529 ( .Z(N6107), .A(N4), .B(N5462) );
and4_1 U1530 ( .Z(N6108), .A(N5549), .B(N5488), .C(N5477), .D(N5470) );
and2_1 U1531 ( .Z(N6111), .A(N5477), .B(N4320) );
and3_1 U1532 ( .Z(N6112), .A(N5488), .B(N4325), .C(N5477) );
and3_1 U1533 ( .Z(N6113), .A(N5549), .B(N5488), .C(N5477) );
and2_1 U1534 ( .Z(N6114), .A(N5477), .B(N4320) );
and3_1 U1535 ( .Z(N6115), .A(N5488), .B(N4325), .C(N5477) );
and2_1 U1536 ( .Z(N6116), .A(N5488), .B(N4325) );
and5_1 U1537 ( .Z(N6117), .A(N5555), .B(N5536), .C(N5520), .D(N5506), .E(N5498) );
and2_1 U1538 ( .Z(N6120), .A(N5498), .B(N4332) );
and3_1 U1539 ( .Z(N6121), .A(N5506), .B(N5498), .C(N4336) );
and4_1 U1540 ( .Z(N6122), .A(N5520), .B(N5498), .C(N4342), .D(N5506) );
and5_1 U1541 ( .Z(N6123), .A(N5536), .B(N5520), .C(N5498), .D(N4349), .E(N5506) );
and2_1 U1542 ( .Z(N6124), .A(N5506), .B(N4336) );
and3_1 U1543 ( .Z(N6125), .A(N5520), .B(N4342), .C(N5506) );
and4_1 U1544 ( .Z(N6126), .A(N5536), .B(N5520), .C(N4349), .D(N5506) );
and4_1 U1545 ( .Z(N6127), .A(N5555), .B(N5520), .C(N5506), .D(N5536) );
and2_1 U1546 ( .Z(N6128), .A(N5506), .B(N4336) );
and3_1 U1547 ( .Z(N6129), .A(N5520), .B(N4342), .C(N5506) );
and4_1 U1548 ( .Z(N6130), .A(N5536), .B(N5520), .C(N4349), .D(N5506) );
and2_1 U1549 ( .Z(N6131), .A(N5520), .B(N4342) );
and3_1 U1550 ( .Z(N6132), .A(N5536), .B(N5520), .C(N4349) );
and3_1 U1551 ( .Z(N6133), .A(N5555), .B(N5520), .C(N5536) );
and2_1 U1552 ( .Z(N6134), .A(N5520), .B(N4342) );
and3_1 U1553 ( .Z(N6135), .A(N5536), .B(N5520), .C(N4349) );
and2_1 U1554 ( .Z(N6136), .A(N5536), .B(N4349) );
and2_1 U1555 ( .Z(N6137), .A(N5549), .B(N5488) );
and2_1 U1556 ( .Z(N6138), .A(N5555), .B(N5536) );
inv_1 U1557 ( .Z(N6139), .A(N5573) );
and4_1 U1558 ( .Z(N6140), .A(N4364), .B(N5573), .C(N5562), .D(N4357) );
and3_1 U1559 ( .Z(N6143), .A(N5562), .B(N4385), .C(N4364) );
and3_1 U1560 ( .Z(N6144), .A(N5573), .B(N5562), .C(N4364) );
and3_1 U1561 ( .Z(N6145), .A(N4385), .B(N5562), .C(N4364) );
and2_1 U1562 ( .Z(N6146), .A(N5562), .B(N4385) );
and2_1 U1563 ( .Z(N6147), .A(N5573), .B(N5562) );
and2_1 U1564 ( .Z(N6148), .A(N5562), .B(N4385) );
and5_1 U1565 ( .Z(N6149), .A(N5264), .B(N4405), .C(N5595), .D(N5579), .E(N5606) );
and2_1 U1566 ( .Z(N6152), .A(N5579), .B(N4067) );
and3_1 U1567 ( .Z(N6153), .A(N5264), .B(N5579), .C(N4396) );
and4_1 U1568 ( .Z(N6154), .A(N5595), .B(N5579), .C(N4400), .D(N5264) );
and5_1 U1569 ( .Z(N6155), .A(N5606), .B(N5595), .C(N5579), .D(N4412), .E(N5264) );
and3_1 U1570 ( .Z(N6156), .A(N5595), .B(N4400), .C(N5264) );
and4_1 U1571 ( .Z(N6157), .A(N5606), .B(N5595), .C(N4412), .D(N5264) );
and5_1 U1572 ( .Z(N6158), .A(N54), .B(N4405), .C(N5595), .D(N5606), .E(N5264) );
and2_1 U1573 ( .Z(N6159), .A(N4400), .B(N5595) );
and3_1 U1574 ( .Z(N6160), .A(N5606), .B(N5595), .C(N4412) );
and4_1 U1575 ( .Z(N6161), .A(N54), .B(N4405), .C(N5595), .D(N5606) );
and2_1 U1576 ( .Z(N6162), .A(N5606), .B(N4412) );
and3_1 U1577 ( .Z(N6163), .A(N54), .B(N4405), .C(N5606) );
nand2_1 U1578 ( .Z(N6164), .A(N5616), .B(N5955) );
and4_1 U1579 ( .Z(N6168), .A(N5684), .B(N5624), .C(N4425), .D(N4418) );
and3_1 U1580 ( .Z(N6171), .A(N5624), .B(N4445), .C(N4425) );
and3_1 U1581 ( .Z(N6172), .A(N5684), .B(N5624), .C(N4425) );
and3_1 U1582 ( .Z(N6173), .A(N5624), .B(N4445), .C(N4425) );
and2_1 U1583 ( .Z(N6174), .A(N5624), .B(N4445) );
and5_1 U1584 ( .Z(N6175), .A(N4477), .B(N5671), .C(N5655), .D(N5284), .E(N5634) );
and2_1 U1585 ( .Z(N6178), .A(N5634), .B(N4080) );
and3_1 U1586 ( .Z(N6179), .A(N5284), .B(N5634), .C(N4456) );
and4_1 U1587 ( .Z(N6180), .A(N5655), .B(N5634), .C(N4462), .D(N5284) );
and5_1 U1588 ( .Z(N6181), .A(N5671), .B(N5655), .C(N5634), .D(N4469), .E(N5284) );
and3_1 U1589 ( .Z(N6182), .A(N5655), .B(N4462), .C(N5284) );
and4_1 U1590 ( .Z(N6183), .A(N5671), .B(N5655), .C(N4469), .D(N5284) );
and4_1 U1591 ( .Z(N6184), .A(N4477), .B(N5655), .C(N5284), .D(N5671) );
and3_1 U1592 ( .Z(N6185), .A(N5655), .B(N4462), .C(N5284) );
and4_1 U1593 ( .Z(N6186), .A(N5671), .B(N5655), .C(N4469), .D(N5284) );
and2_1 U1594 ( .Z(N6187), .A(N5655), .B(N4462) );
and3_1 U1595 ( .Z(N6188), .A(N5671), .B(N5655), .C(N4469) );
and3_1 U1596 ( .Z(N6189), .A(N4477), .B(N5655), .C(N5671) );
and2_1 U1597 ( .Z(N6190), .A(N5655), .B(N4462) );
and3_1 U1598 ( .Z(N6191), .A(N5671), .B(N5655), .C(N4469) );
and2_1 U1599 ( .Z(N6192), .A(N5671), .B(N4469) );
and2_1 U1600 ( .Z(N6193), .A(N5684), .B(N5624) );
and2_1 U1601 ( .Z(N6194), .A(N4477), .B(N5671) );
inv_1 U1602 ( .Z(N6197), .A(N5692) );
inv_1 U1603 ( .Z(N6200), .A(N5696) );
inv_1 U1604 ( .Z(N6203), .A(N5703) );
inv_1 U1605 ( .Z(N6206), .A(N5707) );
buf_1 U1606 ( .Z(N6209), .A(N5700) );
buf_1 U1607 ( .Z(N6212), .A(N5700) );
buf_1 U1608 ( .Z(N6215), .A(N5711) );
buf_1 U1609 ( .Z(N6218), .A(N5711) );
nand2_1 U1610 ( .Z(N6221), .A(N5049), .B(N6023) );
inv_1 U1611 ( .Z(N6234), .A(N5756) );
nand2_1 U1612 ( .Z(N6235), .A(N5756), .B(N6044) );
buf_1 U1613 ( .Z(N6238), .A(N5462) );
buf_1 U1614 ( .Z(N6241), .A(N5389) );
buf_1 U1615 ( .Z(N6244), .A(N5389) );
buf_1 U1616 ( .Z(N6247), .A(N5396) );
buf_1 U1617 ( .Z(N6250), .A(N5396) );
buf_1 U1618 ( .Z(N6253), .A(N5407) );
buf_1 U1619 ( .Z(N6256), .A(N5407) );
buf_1 U1620 ( .Z(N6259), .A(N5424) );
buf_1 U1621 ( .Z(N6262), .A(N5431) );
buf_1 U1622 ( .Z(N6265), .A(N5441) );
buf_1 U1623 ( .Z(N6268), .A(N5452) );
buf_1 U1624 ( .Z(N6271), .A(N5549) );
buf_1 U1625 ( .Z(N6274), .A(N5488) );
buf_1 U1626 ( .Z(N6277), .A(N5470) );
buf_1 U1627 ( .Z(N6280), .A(N5477) );
buf_1 U1628 ( .Z(N6283), .A(N5549) );
buf_1 U1629 ( .Z(N6286), .A(N5488) );
buf_1 U1630 ( .Z(N6289), .A(N5470) );
buf_1 U1631 ( .Z(N6292), .A(N5477) );
buf_1 U1632 ( .Z(N6295), .A(N5555) );
buf_1 U1633 ( .Z(N6298), .A(N5536) );
buf_1 U1634 ( .Z(N6301), .A(N5498) );
buf_1 U1635 ( .Z(N6304), .A(N5520) );
buf_1 U1636 ( .Z(N6307), .A(N5506) );
buf_1 U1637 ( .Z(N6310), .A(N5506) );
buf_1 U1638 ( .Z(N6313), .A(N5555) );
buf_1 U1639 ( .Z(N6316), .A(N5536) );
buf_1 U1640 ( .Z(N6319), .A(N5498) );
buf_1 U1641 ( .Z(N6322), .A(N5520) );
buf_1 U1642 ( .Z(N6325), .A(N5562) );
buf_1 U1643 ( .Z(N6328), .A(N5562) );
buf_1 U1644 ( .Z(N6331), .A(N5579) );
buf_1 U1645 ( .Z(N6335), .A(N5595) );
buf_1 U1646 ( .Z(N6338), .A(N5606) );
buf_1 U1647 ( .Z(N6341), .A(N5684) );
buf_1 U1648 ( .Z(N6344), .A(N5624) );
buf_1 U1649 ( .Z(N6347), .A(N5684) );
buf_1 U1650 ( .Z(N6350), .A(N5624) );
buf_1 U1651 ( .Z(N6353), .A(N5671) );
buf_1 U1652 ( .Z(N6356), .A(N5634) );
buf_1 U1653 ( .Z(N6359), .A(N5655) );
buf_1 U1654 ( .Z(N6364), .A(N5671) );
buf_1 U1655 ( .Z(N6367), .A(N5634) );
buf_1 U1656 ( .Z(N6370), .A(N5655) );
inv_1 U1657 ( .Z(N6373), .A(N5736) );
inv_1 U1658 ( .Z(N6374), .A(N5739) );
inv_1 U1659 ( .Z(N6375), .A(N5742) );
inv_1 U1660 ( .Z(N6376), .A(N5745) );
nand2_1 U1661 ( .Z(N6377), .A(N4243), .B(N6065) );
nand2_1 U1662 ( .Z(N6378), .A(N5236), .B(N6068) );
or4_1 U1663 ( .Z(N6382), .A(N4268), .B(N6071), .C(N6072), .D(N6073) );
or4_1 U1664 ( .Z(N6386), .A(N3968), .B(N5065), .C(N5066), .D(N6074) );
or4_1 U1665 ( .Z(N6388), .A(N4271), .B(N6075), .C(N6076), .D(N6077) );
or4_1 U1666 ( .Z(N6392), .A(N3968), .B(N5067), .C(N5068), .D(N6078) );
or5_1 U1667 ( .Z(N6397), .A(N4297), .B(N6094), .C(N6095), .D(N6096), .E(N6097) );
or2_1 U1668 ( .Z(N6411), .A(N4320), .B(N6116) );
or5_1 U1669 ( .Z(N6415), .A(N4331), .B(N6120), .C(N6121), .D(N6122), .E(N6123) );
or2_1 U1670 ( .Z(N6419), .A(N4342), .B(N6136) );
or5_1 U1671 ( .Z(N6427), .A(N4392), .B(N6152), .C(N6153), .D(N6154), .E(N6155) );
inv_1 U1672 ( .Z(N6434), .A(N6048) );
or2_1 U1673 ( .Z(N6437), .A(N4440), .B(N6174) );
or5_1 U1674 ( .Z(N6441), .A(N4451), .B(N6178), .C(N6179), .D(N6180), .E(N6181) );
or2_1 U1675 ( .Z(N6445), .A(N4462), .B(N6192) );
inv_1 U1676 ( .Z(N6448), .A(N6051) );
inv_1 U1677 ( .Z(N6449), .A(N6054) );
nand2_1 U1678 ( .Z(N6466), .A(N6221), .B(N6024) );
inv_1 U1679 ( .Z(N6469), .A(N6031) );
inv_1 U1680 ( .Z(N6470), .A(N6034) );
inv_1 U1681 ( .Z(N6471), .A(N6037) );
inv_1 U1682 ( .Z(N6472), .A(N6040) );
and3_1 U1683 ( .Z(N6473), .A(N5315), .B(N4524), .C(N6031) );
and3_1 U1684 ( .Z(N6474), .A(N6025), .B(N5150), .C(N6034) );
and3_1 U1685 ( .Z(N6475), .A(N5324), .B(N4532), .C(N6037) );
and3_1 U1686 ( .Z(N6476), .A(N6028), .B(N5157), .C(N6040) );
nand2_1 U1687 ( .Z(N6477), .A(N5385), .B(N6234) );
nand2_1 U1688 ( .Z(N6478), .A(N6045), .B(N132) );
or4_1 U1689 ( .Z(N6482), .A(N4280), .B(N6083), .C(N6084), .D(N6085) );
nor3_1 U1690 ( .Z(N6486), .A(N4280), .B(N6086), .C(N6087) );
or3_1 U1691 ( .Z(N6490), .A(N4284), .B(N6088), .C(N6089) );
nor2_1 U1692 ( .Z(N6494), .A(N4284), .B(N6090) );
or5_1 U1693 ( .Z(N6500), .A(N4298), .B(N6098), .C(N6099), .D(N6100), .E(N6101) );
or4_1 U1694 ( .Z(N6504), .A(N4301), .B(N6102), .C(N6103), .D(N6104) );
or3_1 U1695 ( .Z(N6508), .A(N4305), .B(N6105), .C(N6106) );
or2_1 U1696 ( .Z(N6512), .A(N4310), .B(N6107) );
or4_1 U1697 ( .Z(N6516), .A(N4316), .B(N6111), .C(N6112), .D(N6113) );
nor3_1 U1698 ( .Z(N6526), .A(N4316), .B(N6114), .C(N6115) );
or4_1 U1699 ( .Z(N6536), .A(N4336), .B(N6131), .C(N6132), .D(N6133) );
or5_1 U1700 ( .Z(N6539), .A(N4332), .B(N6124), .C(N6125), .D(N6126), .E(N6127) );
nor3_1 U1701 ( .Z(N6553), .A(N4336), .B(N6134), .C(N6135) );
nor4_1 U1702 ( .Z(N6556), .A(N4332), .B(N6128), .C(N6129), .D(N6130) );
or4_1 U1703 ( .Z(N6566), .A(N4375), .B(N5117), .C(N6143), .D(N6144) );
nor3_1 U1704 ( .Z(N6569), .A(N4375), .B(N5118), .C(N6145) );
or3_1 U1705 ( .Z(N6572), .A(N4379), .B(N6146), .C(N6147) );
nor2_1 U1706 ( .Z(N6575), .A(N4379), .B(N6148) );
or5_1 U1707 ( .Z(N6580), .A(N4067), .B(N5954), .C(N6156), .D(N6157), .E(N6158) );
or4_1 U1708 ( .Z(N6584), .A(N4396), .B(N6159), .C(N6160), .D(N6161) );
or3_1 U1709 ( .Z(N6587), .A(N4400), .B(N6162), .C(N6163) );
or4_1 U1710 ( .Z(N6592), .A(N4436), .B(N5132), .C(N6171), .D(N6172) );
nor3_1 U1711 ( .Z(N6599), .A(N4436), .B(N5133), .C(N6173) );
or4_1 U1712 ( .Z(N6606), .A(N4456), .B(N6187), .C(N6188), .D(N6189) );
or5_1 U1713 ( .Z(N6609), .A(N4080), .B(N6005), .C(N6182), .D(N6183), .E(N6184) );
nor3_1 U1714 ( .Z(N6619), .A(N4456), .B(N6190), .C(N6191) );
nor4_1 U1715 ( .Z(N6622), .A(N4080), .B(N6006), .C(N6185), .D(N6186) );
nand2_1 U1716 ( .Z(N6630), .A(N5739), .B(N6373) );
nand2_1 U1717 ( .Z(N6631), .A(N5736), .B(N6374) );
nand2_1 U1718 ( .Z(N6632), .A(N5745), .B(N6375) );
nand2_1 U1719 ( .Z(N6633), .A(N5742), .B(N6376) );
nand2_1 U1720 ( .Z(N6634), .A(N6377), .B(N6066) );
nand2_1 U1721 ( .Z(N6637), .A(N6069), .B(N6378) );
inv_1 U1722 ( .Z(N6640), .A(N6164) );
and2_1 U1723 ( .Z(N6641), .A(N6108), .B(N6117) );
and2_1 U1724 ( .Z(N6643), .A(N6140), .B(N6149) );
and2_1 U1725 ( .Z(N6646), .A(N6168), .B(N6175) );
and2_1 U1726 ( .Z(N6648), .A(N6080), .B(N6091) );
nand2_1 U1727 ( .Z(N6650), .A(N6238), .B(N2637) );
inv_1 U1728 ( .Z(N6651), .A(N6238) );
inv_1 U1729 ( .Z(N6653), .A(N6241) );
inv_1 U1730 ( .Z(N6655), .A(N6244) );
inv_1 U1731 ( .Z(N6657), .A(N6247) );
inv_1 U1732 ( .Z(N6659), .A(N6250) );
nand2_1 U1733 ( .Z(N6660), .A(N6253), .B(N5087) );
inv_1 U1734 ( .Z(N6661), .A(N6253) );
nand2_1 U1735 ( .Z(N6662), .A(N6256), .B(N5469) );
inv_1 U1736 ( .Z(N6663), .A(N6256) );
and2_1 U1737 ( .Z(N6664), .A(N6091), .B(N4) );
inv_1 U1738 ( .Z(N6666), .A(N6259) );
inv_1 U1739 ( .Z(N6668), .A(N6262) );
inv_1 U1740 ( .Z(N6670), .A(N6265) );
inv_1 U1741 ( .Z(N6672), .A(N6268) );
inv_1 U1742 ( .Z(N6675), .A(N6117) );
inv_1 U1743 ( .Z(N6680), .A(N6280) );
inv_1 U1744 ( .Z(N6681), .A(N6292) );
inv_1 U1745 ( .Z(N6682), .A(N6307) );
inv_1 U1746 ( .Z(N6683), .A(N6310) );
nand2_1 U1747 ( .Z(N6689), .A(N6325), .B(N5120) );
inv_1 U1748 ( .Z(N6690), .A(N6325) );
nand2_1 U1749 ( .Z(N6691), .A(N6328), .B(N5622) );
inv_1 U1750 ( .Z(N6692), .A(N6328) );
and2_1 U1751 ( .Z(N6693), .A(N6149), .B(N54) );
inv_1 U1752 ( .Z(N6695), .A(N6331) );
inv_1 U1753 ( .Z(N6698), .A(N6335) );
nand2_1 U1754 ( .Z(N6699), .A(N6338), .B(N5956) );
inv_1 U1755 ( .Z(N6700), .A(N6338) );
inv_1 U1756 ( .Z(N6703), .A(N6175) );
inv_1 U1757 ( .Z(N6708), .A(N6209) );
inv_1 U1758 ( .Z(N6709), .A(N6212) );
inv_1 U1759 ( .Z(N6710), .A(N6215) );
inv_1 U1760 ( .Z(N6711), .A(N6218) );
and3_1 U1761 ( .Z(N6712), .A(N5696), .B(N5692), .C(N6209) );
and3_1 U1762 ( .Z(N6713), .A(N6200), .B(N6197), .C(N6212) );
and3_1 U1763 ( .Z(N6714), .A(N5707), .B(N5703), .C(N6215) );
and3_1 U1764 ( .Z(N6715), .A(N6206), .B(N6203), .C(N6218) );
buf_1 U1765 ( .Z(N6716), .A(N6466) );
and3_1 U1766 ( .Z(N6718), .A(N6164), .B(N1777), .C(N3130) );
and3_1 U1767 ( .Z(N6719), .A(N5150), .B(N5315), .C(N6469) );
and3_1 U1768 ( .Z(N6720), .A(N4524), .B(N6025), .C(N6470) );
and3_1 U1769 ( .Z(N6721), .A(N5157), .B(N5324), .C(N6471) );
and3_1 U1770 ( .Z(N6722), .A(N4532), .B(N6028), .C(N6472) );
nand2_1 U1771 ( .Z(N6724), .A(N6477), .B(N6235) );
inv_1 U1772 ( .Z(N6739), .A(N6271) );
inv_1 U1773 ( .Z(N6740), .A(N6274) );
inv_1 U1774 ( .Z(N6741), .A(N6277) );
inv_1 U1775 ( .Z(N6744), .A(N6283) );
inv_1 U1776 ( .Z(N6745), .A(N6286) );
inv_1 U1777 ( .Z(N6746), .A(N6289) );
inv_1 U1778 ( .Z(N6751), .A(N6295) );
inv_1 U1779 ( .Z(N6752), .A(N6298) );
inv_1 U1780 ( .Z(N6753), .A(N6301) );
inv_1 U1781 ( .Z(N6754), .A(N6304) );
inv_1 U1782 ( .Z(N6755), .A(N6322) );
inv_1 U1783 ( .Z(N6760), .A(N6313) );
inv_1 U1784 ( .Z(N6761), .A(N6316) );
inv_1 U1785 ( .Z(N6762), .A(N6319) );
inv_1 U1786 ( .Z(N6772), .A(N6341) );
inv_1 U1787 ( .Z(N6773), .A(N6344) );
inv_1 U1788 ( .Z(N6776), .A(N6347) );
inv_1 U1789 ( .Z(N6777), .A(N6350) );
inv_1 U1790 ( .Z(N6782), .A(N6353) );
inv_1 U1791 ( .Z(N6783), .A(N6356) );
inv_1 U1792 ( .Z(N6784), .A(N6359) );
inv_1 U1793 ( .Z(N6785), .A(N6370) );
inv_1 U1794 ( .Z(N6790), .A(N6364) );
inv_1 U1795 ( .Z(N6791), .A(N6367) );
nand2_1 U1796 ( .Z(N6792), .A(N6630), .B(N6631) );
nand2_1 U1797 ( .Z(N6795), .A(N6632), .B(N6633) );
and2_1 U1798 ( .Z(N6801), .A(N6108), .B(N6415) );
and2_1 U1799 ( .Z(N6802), .A(N6427), .B(N6140) );
and2_1 U1800 ( .Z(N6803), .A(N6397), .B(N6080) );
and2_1 U1801 ( .Z(N6804), .A(N6168), .B(N6441) );
inv_1 U1802 ( .Z(N6805), .A(N6466) );
nand2_1 U1803 ( .Z(N6806), .A(N1851), .B(N6651) );
inv_1 U1804 ( .Z(N6807), .A(N6482) );
nand2_1 U1805 ( .Z(N6808), .A(N6482), .B(N6653) );
inv_1 U1806 ( .Z(N6809), .A(N6486) );
nand2_1 U1807 ( .Z(N6810), .A(N6486), .B(N6655) );
inv_1 U1808 ( .Z(N6811), .A(N6490) );
nand2_1 U1809 ( .Z(N6812), .A(N6490), .B(N6657) );
inv_1 U1810 ( .Z(N6813), .A(N6494) );
nand2_1 U1811 ( .Z(N6814), .A(N6494), .B(N6659) );
nand2_1 U1812 ( .Z(N6815), .A(N4575), .B(N6661) );
nand2_1 U1813 ( .Z(N6816), .A(N5169), .B(N6663) );
or2_1 U1814 ( .Z(N6817), .A(N6397), .B(N6664) );
inv_1 U1815 ( .Z(N6823), .A(N6500) );
nand2_1 U1816 ( .Z(N6824), .A(N6500), .B(N6666) );
inv_1 U1817 ( .Z(N6825), .A(N6504) );
nand2_1 U1818 ( .Z(N6826), .A(N6504), .B(N6668) );
inv_1 U1819 ( .Z(N6827), .A(N6508) );
nand2_1 U1820 ( .Z(N6828), .A(N6508), .B(N6670) );
inv_1 U1821 ( .Z(N6829), .A(N6512) );
nand2_1 U1822 ( .Z(N6830), .A(N6512), .B(N6672) );
inv_1 U1823 ( .Z(N6831), .A(N6415) );
inv_1 U1824 ( .Z(N6834), .A(N6566) );
nand2_1 U1825 ( .Z(N6835), .A(N6566), .B(N5618) );
inv_1 U1826 ( .Z(N6836), .A(N6569) );
nand2_1 U1827 ( .Z(N6837), .A(N6569), .B(N5619) );
inv_1 U1828 ( .Z(N6838), .A(N6572) );
nand2_1 U1829 ( .Z(N6839), .A(N6572), .B(N5620) );
inv_1 U1830 ( .Z(N6840), .A(N6575) );
nand2_1 U1831 ( .Z(N6841), .A(N6575), .B(N5621) );
nand2_1 U1832 ( .Z(N6842), .A(N4627), .B(N6690) );
nand2_1 U1833 ( .Z(N6843), .A(N5195), .B(N6692) );
or2_1 U1834 ( .Z(N6844), .A(N6427), .B(N6693) );
inv_1 U1835 ( .Z(N6850), .A(N6580) );
nand2_1 U1836 ( .Z(N6851), .A(N6580), .B(N6695) );
inv_1 U1837 ( .Z(N6852), .A(N6584) );
nand2_1 U1838 ( .Z(N6853), .A(N6584), .B(N6434) );
inv_1 U1839 ( .Z(N6854), .A(N6587) );
nand2_1 U1840 ( .Z(N6855), .A(N6587), .B(N6698) );
nand2_1 U1841 ( .Z(N6856), .A(N5346), .B(N6700) );
inv_1 U1842 ( .Z(N6857), .A(N6441) );
and3_1 U1843 ( .Z(N6860), .A(N6197), .B(N5696), .C(N6708) );
and3_1 U1844 ( .Z(N6861), .A(N5692), .B(N6200), .C(N6709) );
and3_1 U1845 ( .Z(N6862), .A(N6203), .B(N5707), .C(N6710) );
and3_1 U1846 ( .Z(N6863), .A(N5703), .B(N6206), .C(N6711) );
or3_1 U1847 ( .Z(N6866), .A(N4197), .B(N6718), .C(N3785) );
nor2_1 U1848 ( .Z(N6872), .A(N6719), .B(N6473) );
nor2_1 U1849 ( .Z(N6873), .A(N6720), .B(N6474) );
nor2_1 U1850 ( .Z(N6874), .A(N6721), .B(N6475) );
nor2_1 U1851 ( .Z(N6875), .A(N6722), .B(N6476) );
inv_1 U1852 ( .Z(N6876), .A(N6637) );
buf_1 U1853 ( .Z(N6877), .A(N6724) );
and2_1 U1854 ( .Z(N6879), .A(N6045), .B(N6478) );
and2_1 U1855 ( .Z(N6880), .A(N6478), .B(N132) );
or2_1 U1856 ( .Z(N6881), .A(N6411), .B(N6137) );
inv_1 U1857 ( .Z(N6884), .A(N6516) );
inv_1 U1858 ( .Z(N6885), .A(N6411) );
inv_1 U1859 ( .Z(N6888), .A(N6526) );
inv_1 U1860 ( .Z(N6889), .A(N6536) );
nand2_1 U1861 ( .Z(N6890), .A(N6536), .B(N5176) );
or2_1 U1862 ( .Z(N6891), .A(N6419), .B(N6138) );
inv_1 U1863 ( .Z(N6894), .A(N6539) );
inv_1 U1864 ( .Z(N6895), .A(N6553) );
nand2_1 U1865 ( .Z(N6896), .A(N6553), .B(N5728) );
inv_1 U1866 ( .Z(N6897), .A(N6419) );
inv_1 U1867 ( .Z(N6900), .A(N6556) );
or2_1 U1868 ( .Z(N6901), .A(N6437), .B(N6193) );
inv_1 U1869 ( .Z(N6904), .A(N6592) );
inv_1 U1870 ( .Z(N6905), .A(N6437) );
inv_1 U1871 ( .Z(N6908), .A(N6599) );
or2_1 U1872 ( .Z(N6909), .A(N6445), .B(N6194) );
inv_1 U1873 ( .Z(N6912), .A(N6606) );
inv_1 U1874 ( .Z(N6913), .A(N6609) );
inv_1 U1875 ( .Z(N6914), .A(N6619) );
nand2_1 U1876 ( .Z(N6915), .A(N6619), .B(N5734) );
inv_1 U1877 ( .Z(N6916), .A(N6445) );
inv_1 U1878 ( .Z(N6919), .A(N6622) );
inv_1 U1879 ( .Z(N6922), .A(N6634) );
nand2_1 U1880 ( .Z(N6923), .A(N6634), .B(N6067) );
or2_1 U1881 ( .Z(N6924), .A(N6382), .B(N6801) );
or2_1 U1882 ( .Z(N6925), .A(N6386), .B(N6802) );
or2_1 U1883 ( .Z(N6926), .A(N6388), .B(N6803) );
or2_1 U1884 ( .Z(N6927), .A(N6392), .B(N6804) );
inv_1 U1885 ( .Z(N6930), .A(N6724) );
nand2_1 U1886 ( .Z(N6932), .A(N6650), .B(N6806) );
nand2_1 U1887 ( .Z(N6935), .A(N6241), .B(N6807) );
nand2_1 U1888 ( .Z(N6936), .A(N6244), .B(N6809) );
nand2_1 U1889 ( .Z(N6937), .A(N6247), .B(N6811) );
nand2_1 U1890 ( .Z(N6938), .A(N6250), .B(N6813) );
nand2_1 U1891 ( .Z(N6939), .A(N6660), .B(N6815) );
nand2_1 U1892 ( .Z(N6940), .A(N6662), .B(N6816) );
nand2_1 U1893 ( .Z(N6946), .A(N6259), .B(N6823) );
nand2_1 U1894 ( .Z(N6947), .A(N6262), .B(N6825) );
nand2_1 U1895 ( .Z(N6948), .A(N6265), .B(N6827) );
nand2_1 U1896 ( .Z(N6949), .A(N6268), .B(N6829) );
nand2_1 U1897 ( .Z(N6953), .A(N5183), .B(N6834) );
nand2_1 U1898 ( .Z(N6954), .A(N5186), .B(N6836) );
nand2_1 U1899 ( .Z(N6955), .A(N5189), .B(N6838) );
nand2_1 U1900 ( .Z(N6956), .A(N5192), .B(N6840) );
nand2_1 U1901 ( .Z(N6957), .A(N6689), .B(N6842) );
nand2_1 U1902 ( .Z(N6958), .A(N6691), .B(N6843) );
nand2_1 U1903 ( .Z(N6964), .A(N6331), .B(N6850) );
nand2_1 U1904 ( .Z(N6965), .A(N6048), .B(N6852) );
nand2_1 U1905 ( .Z(N6966), .A(N6335), .B(N6854) );
nand2_1 U1906 ( .Z(N6967), .A(N6699), .B(N6856) );
nor2_1 U1907 ( .Z(N6973), .A(N6860), .B(N6712) );
nor2_1 U1908 ( .Z(N6974), .A(N6861), .B(N6713) );
nor2_1 U1909 ( .Z(N6975), .A(N6862), .B(N6714) );
nor2_1 U1910 ( .Z(N6976), .A(N6863), .B(N6715) );
inv_1 U1911 ( .Z(N6977), .A(N6792) );
inv_1 U1912 ( .Z(N6978), .A(N6795) );
or2_1 U1913 ( .Z(N6979), .A(N6879), .B(N6880) );
nand2_1 U1914 ( .Z(N6987), .A(N4608), .B(N6889) );
nand2_1 U1915 ( .Z(N6990), .A(N5177), .B(N6895) );
nand2_1 U1916 ( .Z(N6999), .A(N5217), .B(N6914) );
nand2_1 U1917 ( .Z(N7002), .A(N5377), .B(N6922) );
nand2_1 U1918 ( .Z(N7003), .A(N6873), .B(N6872) );
nand2_1 U1919 ( .Z(N7006), .A(N6875), .B(N6874) );
and3_1 U1920 ( .Z(N7011), .A(N6866), .B(N2681), .C(N2692) );
and3_1 U1921 ( .Z(N7012), .A(N6866), .B(N2756), .C(N2767) );
and3_1 U1922 ( .Z(N7013), .A(N6866), .B(N2779), .C(N2790) );
inv_1 U1923 ( .Z(N7015), .A(N6866) );
and3_1 U1924 ( .Z(N7016), .A(N6866), .B(N2801), .C(N2812) );
nand2_1 U1925 ( .Z(N7018), .A(N6935), .B(N6808) );
nand2_1 U1926 ( .Z(N7019), .A(N6936), .B(N6810) );
nand2_1 U1927 ( .Z(N7020), .A(N6937), .B(N6812) );
nand2_1 U1928 ( .Z(N7021), .A(N6938), .B(N6814) );
inv_1 U1929 ( .Z(N7022), .A(N6939) );
inv_1 U1930 ( .Z(N7023), .A(N6817) );
nand2_1 U1931 ( .Z(N7028), .A(N6946), .B(N6824) );
nand2_1 U1932 ( .Z(N7031), .A(N6947), .B(N6826) );
nand2_1 U1933 ( .Z(N7034), .A(N6948), .B(N6828) );
nand2_1 U1934 ( .Z(N7037), .A(N6949), .B(N6830) );
and2_1 U1935 ( .Z(N7040), .A(N6817), .B(N6079) );
and2_1 U1936 ( .Z(N7041), .A(N6831), .B(N6675) );
nand2_1 U1937 ( .Z(N7044), .A(N6953), .B(N6835) );
nand2_1 U1938 ( .Z(N7045), .A(N6954), .B(N6837) );
nand2_1 U1939 ( .Z(N7046), .A(N6955), .B(N6839) );
nand2_1 U1940 ( .Z(N7047), .A(N6956), .B(N6841) );
inv_1 U1941 ( .Z(N7048), .A(N6957) );
inv_1 U1942 ( .Z(N7049), .A(N6844) );
nand2_1 U1943 ( .Z(N7054), .A(N6964), .B(N6851) );
nand2_1 U1944 ( .Z(N7057), .A(N6965), .B(N6853) );
nand2_1 U1945 ( .Z(N7060), .A(N6966), .B(N6855) );
and2_1 U1946 ( .Z(N7064), .A(N6844), .B(N6139) );
and2_1 U1947 ( .Z(N7065), .A(N6857), .B(N6703) );
inv_1 U1948 ( .Z(N7072), .A(N6881) );
nand2_1 U1949 ( .Z(N7073), .A(N6881), .B(N5172) );
inv_1 U1950 ( .Z(N7074), .A(N6885) );
nand2_1 U1951 ( .Z(N7075), .A(N6885), .B(N5727) );
nand2_1 U1952 ( .Z(N7076), .A(N6890), .B(N6987) );
inv_1 U1953 ( .Z(N7079), .A(N6891) );
nand2_1 U1954 ( .Z(N7080), .A(N6896), .B(N6990) );
inv_1 U1955 ( .Z(N7083), .A(N6897) );
inv_1 U1956 ( .Z(N7084), .A(N6901) );
nand2_1 U1957 ( .Z(N7085), .A(N6901), .B(N5198) );
inv_1 U1958 ( .Z(N7086), .A(N6905) );
nand2_1 U1959 ( .Z(N7087), .A(N6905), .B(N5731) );
inv_1 U1960 ( .Z(N7088), .A(N6909) );
nand2_1 U1961 ( .Z(N7089), .A(N6909), .B(N6912) );
nand2_1 U1962 ( .Z(N7090), .A(N6915), .B(N6999) );
inv_1 U1963 ( .Z(N7093), .A(N6916) );
nand2_1 U1964 ( .Z(N7094), .A(N6974), .B(N6973) );
nand2_1 U1965 ( .Z(N7097), .A(N6976), .B(N6975) );
nand2_1 U1966 ( .Z(N7101), .A(N7002), .B(N6923) );
inv_1 U1967 ( .Z(N7105), .A(N6932) );
inv_1 U1968 ( .Z(N7110), .A(N6967) );
and3_1 U1969 ( .Z(N7114), .A(N6979), .B(N603), .C(N1755) );
inv_1 U1970 ( .Z(N7115), .A(N7019) );
inv_1 U1971 ( .Z(N7116), .A(N7021) );
and2_1 U1972 ( .Z(N7125), .A(N6817), .B(N7018) );
and2_1 U1973 ( .Z(N7126), .A(N6817), .B(N7020) );
and2_1 U1974 ( .Z(N7127), .A(N6817), .B(N7022) );
inv_1 U1975 ( .Z(N7130), .A(N7045) );
inv_1 U1976 ( .Z(N7131), .A(N7047) );
and2_1 U1977 ( .Z(N7139), .A(N6844), .B(N7044) );
and2_1 U1978 ( .Z(N7140), .A(N6844), .B(N7046) );
and2_1 U1979 ( .Z(N7141), .A(N6844), .B(N7048) );
and3_1 U1980 ( .Z(N7146), .A(N6932), .B(N1761), .C(N3108) );
and3_1 U1981 ( .Z(N7147), .A(N6967), .B(N1777), .C(N3130) );
inv_1 U1982 ( .Z(N7149), .A(N7003) );
inv_1 U1983 ( .Z(N7150), .A(N7006) );
nand2_1 U1984 ( .Z(N7151), .A(N7006), .B(N6876) );
nand2_1 U1985 ( .Z(N7152), .A(N4605), .B(N7072) );
nand2_1 U1986 ( .Z(N7153), .A(N5173), .B(N7074) );
nand2_1 U1987 ( .Z(N7158), .A(N4646), .B(N7084) );
nand2_1 U1988 ( .Z(N7159), .A(N5205), .B(N7086) );
nand2_1 U1989 ( .Z(N7160), .A(N6606), .B(N7088) );
inv_1 U1990 ( .Z(N7166), .A(N7037) );
inv_1 U1991 ( .Z(N7167), .A(N7034) );
inv_1 U1992 ( .Z(N7168), .A(N7031) );
inv_1 U1993 ( .Z(N7169), .A(N7028) );
inv_1 U1994 ( .Z(N7170), .A(N7060) );
inv_1 U1995 ( .Z(N7171), .A(N7057) );
inv_1 U1996 ( .Z(N7172), .A(N7054) );
and2_1 U1997 ( .Z(N7173), .A(N7115), .B(N7023) );
and2_1 U1998 ( .Z(N7174), .A(N7116), .B(N7023) );
and2_1 U1999 ( .Z(N7175), .A(N6940), .B(N7023) );
and2_1 U2000 ( .Z(N7176), .A(N5418), .B(N7023) );
inv_1 U2001 ( .Z(N7177), .A(N7041) );
and2_1 U2002 ( .Z(N7178), .A(N7130), .B(N7049) );
and2_1 U2003 ( .Z(N7179), .A(N7131), .B(N7049) );
and2_1 U2004 ( .Z(N7180), .A(N6958), .B(N7049) );
and2_1 U2005 ( .Z(N7181), .A(N5573), .B(N7049) );
inv_1 U2006 ( .Z(N7182), .A(N7065) );
inv_1 U2007 ( .Z(N7183), .A(N7094) );
nand2_1 U2008 ( .Z(N7184), .A(N7094), .B(N6977) );
inv_1 U2009 ( .Z(N7185), .A(N7097) );
nand2_1 U2010 ( .Z(N7186), .A(N7097), .B(N6978) );
and3_1 U2011 ( .Z(N7187), .A(N7037), .B(N1761), .C(N3108) );
and3_1 U2012 ( .Z(N7188), .A(N7034), .B(N1761), .C(N3108) );
and3_1 U2013 ( .Z(N7189), .A(N7031), .B(N1761), .C(N3108) );
or3_1 U2014 ( .Z(N7190), .A(N4956), .B(N7146), .C(N3781) );
and3_1 U2015 ( .Z(N7196), .A(N7060), .B(N1777), .C(N3130) );
and3_1 U2016 ( .Z(N7197), .A(N7057), .B(N1777), .C(N3130) );
or3_1 U2017 ( .Z(N7198), .A(N4960), .B(N7147), .C(N3786) );
nand2_1 U2018 ( .Z(N7204), .A(N7101), .B(N7149) );
inv_1 U2019 ( .Z(N7205), .A(N7101) );
nand2_1 U2020 ( .Z(N7206), .A(N6637), .B(N7150) );
and3_1 U2021 ( .Z(N7207), .A(N7028), .B(N1793), .C(N3158) );
and3_1 U2022 ( .Z(N7208), .A(N7054), .B(N1807), .C(N3180) );
nand2_1 U2023 ( .Z(N7209), .A(N7073), .B(N7152) );
nand2_1 U2024 ( .Z(N7212), .A(N7075), .B(N7153) );
inv_1 U2025 ( .Z(N7215), .A(N7076) );
nand2_1 U2026 ( .Z(N7216), .A(N7076), .B(N7079) );
inv_1 U2027 ( .Z(N7217), .A(N7080) );
nand2_1 U2028 ( .Z(N7218), .A(N7080), .B(N7083) );
nand2_1 U2029 ( .Z(N7219), .A(N7085), .B(N7158) );
nand2_1 U2030 ( .Z(N7222), .A(N7087), .B(N7159) );
nand2_1 U2031 ( .Z(N7225), .A(N7089), .B(N7160) );
inv_1 U2032 ( .Z(N7228), .A(N7090) );
nand2_1 U2033 ( .Z(N7229), .A(N7090), .B(N7093) );
or2_1 U2034 ( .Z(N7236), .A(N7173), .B(N7125) );
or2_1 U2035 ( .Z(N7239), .A(N7174), .B(N7126) );
or2_1 U2036 ( .Z(N7242), .A(N7175), .B(N7127) );
or2_1 U2037 ( .Z(N7245), .A(N7176), .B(N7040) );
or2_1 U2038 ( .Z(N7250), .A(N7178), .B(N7139) );
or2_1 U2039 ( .Z(N7257), .A(N7179), .B(N7140) );
or2_1 U2040 ( .Z(N7260), .A(N7180), .B(N7141) );
or2_1 U2041 ( .Z(N7263), .A(N7181), .B(N7064) );
nand2_1 U2042 ( .Z(N7268), .A(N6792), .B(N7183) );
nand2_1 U2043 ( .Z(N7269), .A(N6795), .B(N7185) );
or3_1 U2044 ( .Z(N7270), .A(N4957), .B(N7187), .C(N3782) );
or3_1 U2045 ( .Z(N7276), .A(N4958), .B(N7188), .C(N3783) );
or3_1 U2046 ( .Z(N7282), .A(N4959), .B(N7189), .C(N3784) );
or3_1 U2047 ( .Z(N7288), .A(N4961), .B(N7196), .C(N3787) );
or3_1 U2048 ( .Z(N7294), .A(N3998), .B(N7197), .C(N3788) );
nand2_1 U2049 ( .Z(N7300), .A(N7003), .B(N7205) );
nand2_1 U2050 ( .Z(N7301), .A(N7206), .B(N7151) );
or3_1 U2051 ( .Z(N7304), .A(N4980), .B(N7207), .C(N3800) );
or3_1 U2052 ( .Z(N7310), .A(N4984), .B(N7208), .C(N3805) );
nand2_1 U2053 ( .Z(N7320), .A(N6891), .B(N7215) );
nand2_1 U2054 ( .Z(N7321), .A(N6897), .B(N7217) );
nand2_1 U2055 ( .Z(N7328), .A(N6916), .B(N7228) );
and3_1 U2056 ( .Z(N7338), .A(N7190), .B(N1185), .C(N2692) );
and3_1 U2057 ( .Z(N7339), .A(N7198), .B(N2681), .C(N2692) );
and3_1 U2058 ( .Z(N7340), .A(N7190), .B(N1247), .C(N2767) );
and3_1 U2059 ( .Z(N7341), .A(N7198), .B(N2756), .C(N2767) );
and3_1 U2060 ( .Z(N7342), .A(N7190), .B(N1327), .C(N2790) );
and3_1 U2061 ( .Z(N7349), .A(N7198), .B(N2779), .C(N2790) );
and3_1 U2062 ( .Z(N7357), .A(N7198), .B(N2801), .C(N2812) );
inv_1 U2063 ( .Z(N7363), .A(N7198) );
and3_1 U2064 ( .Z(N7364), .A(N7190), .B(N1351), .C(N2812) );
inv_1 U2065 ( .Z(N7365), .A(N7190) );
nand2_1 U2066 ( .Z(N7394), .A(N7268), .B(N7184) );
nand2_1 U2067 ( .Z(N7397), .A(N7269), .B(N7186) );
nand2_1 U2068 ( .Z(N7402), .A(N7204), .B(N7300) );
inv_1 U2069 ( .Z(N7405), .A(N7209) );
nand2_1 U2070 ( .Z(N7406), .A(N7209), .B(N6884) );
inv_1 U2071 ( .Z(N7407), .A(N7212) );
nand2_1 U2072 ( .Z(N7408), .A(N7212), .B(N6888) );
nand2_1 U2073 ( .Z(N7409), .A(N7320), .B(N7216) );
nand2_1 U2074 ( .Z(N7412), .A(N7321), .B(N7218) );
inv_1 U2075 ( .Z(N7415), .A(N7219) );
nand2_1 U2076 ( .Z(N7416), .A(N7219), .B(N6904) );
inv_1 U2077 ( .Z(N7417), .A(N7222) );
nand2_1 U2078 ( .Z(N7418), .A(N7222), .B(N6908) );
inv_1 U2079 ( .Z(N7419), .A(N7225) );
nand2_1 U2080 ( .Z(N7420), .A(N7225), .B(N6913) );
nand2_1 U2081 ( .Z(N7421), .A(N7328), .B(N7229) );
inv_1 U2082 ( .Z(N7424), .A(N7245) );
inv_1 U2083 ( .Z(N7425), .A(N7242) );
inv_1 U2084 ( .Z(N7426), .A(N7239) );
inv_1 U2085 ( .Z(N7427), .A(N7236) );
inv_1 U2086 ( .Z(N7428), .A(N7263) );
inv_1 U2087 ( .Z(N7429), .A(N7260) );
inv_1 U2088 ( .Z(N7430), .A(N7257) );
inv_1 U2089 ( .Z(N7431), .A(N7250) );
inv_1 U2090 ( .Z(N7432), .A(N7250) );
and3_1 U2091 ( .Z(N7433), .A(N7310), .B(N2653), .C(N2664) );
and3_1 U2092 ( .Z(N7434), .A(N7304), .B(N1161), .C(N2664) );
or4_1 U2093 ( .Z(N7435), .A(N7011), .B(N7338), .C(N3621), .D(N2591) );
and3_1 U2094 ( .Z(N7436), .A(N7270), .B(N1185), .C(N2692) );
and3_1 U2095 ( .Z(N7437), .A(N7288), .B(N2681), .C(N2692) );
and3_1 U2096 ( .Z(N7438), .A(N7276), .B(N1185), .C(N2692) );
and3_1 U2097 ( .Z(N7439), .A(N7294), .B(N2681), .C(N2692) );
and3_1 U2098 ( .Z(N7440), .A(N7282), .B(N1185), .C(N2692) );
and3_1 U2099 ( .Z(N7441), .A(N7310), .B(N2728), .C(N2739) );
and3_1 U2100 ( .Z(N7442), .A(N7304), .B(N1223), .C(N2739) );
or4_1 U2101 ( .Z(N7443), .A(N7012), .B(N7340), .C(N3632), .D(N2600) );
and3_1 U2102 ( .Z(N7444), .A(N7270), .B(N1247), .C(N2767) );
and3_1 U2103 ( .Z(N7445), .A(N7288), .B(N2756), .C(N2767) );
and3_1 U2104 ( .Z(N7446), .A(N7276), .B(N1247), .C(N2767) );
and3_1 U2105 ( .Z(N7447), .A(N7294), .B(N2756), .C(N2767) );
and3_1 U2106 ( .Z(N7448), .A(N7282), .B(N1247), .C(N2767) );
or4_1 U2107 ( .Z(N7449), .A(N7013), .B(N7342), .C(N3641), .D(N2605) );
and3_1 U2108 ( .Z(N7450), .A(N7310), .B(N3041), .C(N3052) );
and3_1 U2109 ( .Z(N7451), .A(N7304), .B(N1697), .C(N3052) );
and3_1 U2110 ( .Z(N7452), .A(N7294), .B(N2779), .C(N2790) );
and3_1 U2111 ( .Z(N7453), .A(N7282), .B(N1327), .C(N2790) );
and3_1 U2112 ( .Z(N7454), .A(N7288), .B(N2779), .C(N2790) );
and3_1 U2113 ( .Z(N7455), .A(N7276), .B(N1327), .C(N2790) );
and3_1 U2114 ( .Z(N7456), .A(N7270), .B(N1327), .C(N2790) );
and3_1 U2115 ( .Z(N7457), .A(N7310), .B(N3075), .C(N3086) );
and3_1 U2116 ( .Z(N7458), .A(N7304), .B(N1731), .C(N3086) );
and3_1 U2117 ( .Z(N7459), .A(N7294), .B(N2801), .C(N2812) );
and3_1 U2118 ( .Z(N7460), .A(N7282), .B(N1351), .C(N2812) );
and3_1 U2119 ( .Z(N7461), .A(N7288), .B(N2801), .C(N2812) );
and3_1 U2120 ( .Z(N7462), .A(N7276), .B(N1351), .C(N2812) );
and3_1 U2121 ( .Z(N7463), .A(N7270), .B(N1351), .C(N2812) );
and3_1 U2122 ( .Z(N7464), .A(N7250), .B(N603), .C(N599) );
inv_1 U2123 ( .Z(N7465), .A(N7310) );
inv_1 U2124 ( .Z(N7466), .A(N7294) );
inv_1 U2125 ( .Z(N7467), .A(N7288) );
inv_1 U2126 ( .Z(N7468), .A(N7301) );
or4_1 U2127 ( .Z(N7469), .A(N7016), .B(N7364), .C(N3660), .D(N2626) );
inv_1 U2128 ( .Z(N7470), .A(N7304) );
inv_1 U2129 ( .Z(N7471), .A(N7282) );
inv_1 U2130 ( .Z(N7472), .A(N7276) );
inv_1 U2131 ( .Z(N7473), .A(N7270) );
buf_1 U2132 ( .Z(N7474), .A(N7394) );
buf_1 U2133 ( .Z(N7476), .A(N7397) );
and2_1 U2134 ( .Z(N7479), .A(N7301), .B(N3068) );
and3_1 U2135 ( .Z(N7481), .A(N7245), .B(N1793), .C(N3158) );
and3_1 U2136 ( .Z(N7482), .A(N7242), .B(N1793), .C(N3158) );
and3_1 U2137 ( .Z(N7483), .A(N7239), .B(N1793), .C(N3158) );
and3_1 U2138 ( .Z(N7484), .A(N7236), .B(N1793), .C(N3158) );
and3_1 U2139 ( .Z(N7485), .A(N7263), .B(N1807), .C(N3180) );
and3_1 U2140 ( .Z(N7486), .A(N7260), .B(N1807), .C(N3180) );
and3_1 U2141 ( .Z(N7487), .A(N7257), .B(N1807), .C(N3180) );
and3_1 U2142 ( .Z(N7488), .A(N7250), .B(N1807), .C(N3180) );
nand2_1 U2143 ( .Z(N7489), .A(N6979), .B(N7250) );
nand2_1 U2144 ( .Z(N7492), .A(N6516), .B(N7405) );
nand2_1 U2145 ( .Z(N7493), .A(N6526), .B(N7407) );
nand2_1 U2146 ( .Z(N7498), .A(N6592), .B(N7415) );
nand2_1 U2147 ( .Z(N7499), .A(N6599), .B(N7417) );
nand2_1 U2148 ( .Z(N7500), .A(N6609), .B(N7419) );
and9_1 U2149 ( .Z(N7503), .A(N7105), .B(N7166), .C(N7167), .D(N7168), .E(N7169), .F(N7424), .G(N7425), .H(N7426), .I(N7427) );
and9_1 U2150 ( .Z(N7504), .A(N6640), .B(N7110), .C(N7170), .D(N7171), .E(N7172), .F(N7428), .G(N7429), .H(N7430), .I(N7431) );
or4_1 U2151 ( .Z(N7505), .A(N7433), .B(N7434), .C(N3616), .D(N2585) );
and2_1 U2152 ( .Z(N7506), .A(N7435), .B(N2675) );
or4_1 U2153 ( .Z(N7507), .A(N7339), .B(N7436), .C(N3622), .D(N2592) );
or4_1 U2154 ( .Z(N7508), .A(N7437), .B(N7438), .C(N3623), .D(N2593) );
or4_1 U2155 ( .Z(N7509), .A(N7439), .B(N7440), .C(N3624), .D(N2594) );
or4_1 U2156 ( .Z(N7510), .A(N7441), .B(N7442), .C(N3627), .D(N2595) );
and2_1 U2157 ( .Z(N7511), .A(N7443), .B(N2750) );
or4_1 U2158 ( .Z(N7512), .A(N7341), .B(N7444), .C(N3633), .D(N2601) );
or4_1 U2159 ( .Z(N7513), .A(N7445), .B(N7446), .C(N3634), .D(N2602) );
or4_1 U2160 ( .Z(N7514), .A(N7447), .B(N7448), .C(N3635), .D(N2603) );
or4_1 U2161 ( .Z(N7515), .A(N7450), .B(N7451), .C(N3646), .D(N2610) );
or4_1 U2162 ( .Z(N7516), .A(N7452), .B(N7453), .C(N3647), .D(N2611) );
or4_1 U2163 ( .Z(N7517), .A(N7454), .B(N7455), .C(N3648), .D(N2612) );
or4_1 U2164 ( .Z(N7518), .A(N7349), .B(N7456), .C(N3649), .D(N2613) );
or4_1 U2165 ( .Z(N7519), .A(N7457), .B(N7458), .C(N3654), .D(N2618) );
or4_1 U2166 ( .Z(N7520), .A(N7459), .B(N7460), .C(N3655), .D(N2619) );
or4_1 U2167 ( .Z(N7521), .A(N7461), .B(N7462), .C(N3656), .D(N2620) );
or4_1 U2168 ( .Z(N7522), .A(N7357), .B(N7463), .C(N3657), .D(N2621) );
or4_1 U2169 ( .Z(N7525), .A(N4741), .B(N7114), .C(N2624), .D(N7464) );
and3_1 U2170 ( .Z(N7526), .A(N7468), .B(N3119), .C(N3130) );
inv_1 U2171 ( .Z(N7527), .A(N7394) );
inv_1 U2172 ( .Z(N7528), .A(N7397) );
inv_1 U2173 ( .Z(N7529), .A(N7402) );
and2_1 U2174 ( .Z(N7530), .A(N7402), .B(N3068) );
or3_1 U2175 ( .Z(N7531), .A(N4981), .B(N7481), .C(N3801) );
or3_1 U2176 ( .Z(N7537), .A(N4982), .B(N7482), .C(N3802) );
or3_1 U2177 ( .Z(N7543), .A(N4983), .B(N7483), .C(N3803) );
or3_1 U2178 ( .Z(N7549), .A(N5165), .B(N7484), .C(N3804) );
or3_1 U2179 ( .Z(N7555), .A(N4985), .B(N7485), .C(N3806) );
or3_1 U2180 ( .Z(N7561), .A(N4986), .B(N7486), .C(N3807) );
or3_1 U2181 ( .Z(N7567), .A(N4547), .B(N7487), .C(N3808) );
or3_1 U2182 ( .Z(N7573), .A(N4987), .B(N7488), .C(N3809) );
nand2_1 U2183 ( .Z(N7579), .A(N7492), .B(N7406) );
nand2_1 U2184 ( .Z(N7582), .A(N7493), .B(N7408) );
inv_1 U2185 ( .Z(N7585), .A(N7409) );
nand2_1 U2186 ( .Z(N7586), .A(N7409), .B(N6894) );
inv_1 U2187 ( .Z(N7587), .A(N7412) );
nand2_1 U2188 ( .Z(N7588), .A(N7412), .B(N6900) );
nand2_1 U2189 ( .Z(N7589), .A(N7498), .B(N7416) );
nand2_1 U2190 ( .Z(N7592), .A(N7499), .B(N7418) );
nand2_1 U2191 ( .Z(N7595), .A(N7500), .B(N7420) );
inv_1 U2192 ( .Z(N7598), .A(N7421) );
nand2_1 U2193 ( .Z(N7599), .A(N7421), .B(N6919) );
and2_1 U2194 ( .Z(N7600), .A(N7505), .B(N2647) );
and2_1 U2195 ( .Z(N7601), .A(N7507), .B(N2675) );
and2_1 U2196 ( .Z(N7602), .A(N7508), .B(N2675) );
and2_1 U2197 ( .Z(N7603), .A(N7509), .B(N2675) );
and2_1 U2198 ( .Z(N7604), .A(N7510), .B(N2722) );
and2_1 U2199 ( .Z(N7605), .A(N7512), .B(N2750) );
and2_1 U2200 ( .Z(N7606), .A(N7513), .B(N2750) );
and2_1 U2201 ( .Z(N7607), .A(N7514), .B(N2750) );
and2_1 U2202 ( .Z(N7624), .A(N6979), .B(N7489) );
and2_1 U2203 ( .Z(N7625), .A(N7489), .B(N7250) );
and2_1 U2204 ( .Z(N7626), .A(N1149), .B(N7525) );
and5_1 U2205 ( .Z(N7631), .A(N562), .B(N7527), .C(N7528), .D(N6805), .E(N6930) );
and3_1 U2206 ( .Z(N7636), .A(N7529), .B(N3097), .C(N3108) );
nand2_1 U2207 ( .Z(N7657), .A(N6539), .B(N7585) );
nand2_1 U2208 ( .Z(N7658), .A(N6556), .B(N7587) );
nand2_1 U2209 ( .Z(N7665), .A(N6622), .B(N7598) );
and3_1 U2210 ( .Z(N7666), .A(N7555), .B(N2653), .C(N2664) );
and3_1 U2211 ( .Z(N7667), .A(N7531), .B(N1161), .C(N2664) );
and3_1 U2212 ( .Z(N7668), .A(N7561), .B(N2653), .C(N2664) );
and3_1 U2213 ( .Z(N7669), .A(N7537), .B(N1161), .C(N2664) );
and3_1 U2214 ( .Z(N7670), .A(N7567), .B(N2653), .C(N2664) );
and3_1 U2215 ( .Z(N7671), .A(N7543), .B(N1161), .C(N2664) );
and3_1 U2216 ( .Z(N7672), .A(N7573), .B(N2653), .C(N2664) );
and3_1 U2217 ( .Z(N7673), .A(N7549), .B(N1161), .C(N2664) );
and3_1 U2218 ( .Z(N7674), .A(N7555), .B(N2728), .C(N2739) );
and3_1 U2219 ( .Z(N7675), .A(N7531), .B(N1223), .C(N2739) );
and3_1 U2220 ( .Z(N7676), .A(N7561), .B(N2728), .C(N2739) );
and3_1 U2221 ( .Z(N7677), .A(N7537), .B(N1223), .C(N2739) );
and3_1 U2222 ( .Z(N7678), .A(N7567), .B(N2728), .C(N2739) );
and3_1 U2223 ( .Z(N7679), .A(N7543), .B(N1223), .C(N2739) );
and3_1 U2224 ( .Z(N7680), .A(N7573), .B(N2728), .C(N2739) );
and3_1 U2225 ( .Z(N7681), .A(N7549), .B(N1223), .C(N2739) );
and3_1 U2226 ( .Z(N7682), .A(N7573), .B(N3075), .C(N3086) );
and3_1 U2227 ( .Z(N7683), .A(N7549), .B(N1731), .C(N3086) );
and3_1 U2228 ( .Z(N7684), .A(N7573), .B(N3041), .C(N3052) );
and3_1 U2229 ( .Z(N7685), .A(N7549), .B(N1697), .C(N3052) );
and3_1 U2230 ( .Z(N7686), .A(N7567), .B(N3041), .C(N3052) );
and3_1 U2231 ( .Z(N7687), .A(N7543), .B(N1697), .C(N3052) );
and3_1 U2232 ( .Z(N7688), .A(N7561), .B(N3041), .C(N3052) );
and3_1 U2233 ( .Z(N7689), .A(N7537), .B(N1697), .C(N3052) );
and3_1 U2234 ( .Z(N7690), .A(N7555), .B(N3041), .C(N3052) );
and3_1 U2235 ( .Z(N7691), .A(N7531), .B(N1697), .C(N3052) );
and3_1 U2236 ( .Z(N7692), .A(N7567), .B(N3075), .C(N3086) );
and3_1 U2237 ( .Z(N7693), .A(N7543), .B(N1731), .C(N3086) );
and3_1 U2238 ( .Z(N7694), .A(N7561), .B(N3075), .C(N3086) );
and3_1 U2239 ( .Z(N7695), .A(N7537), .B(N1731), .C(N3086) );
and3_1 U2240 ( .Z(N7696), .A(N7555), .B(N3075), .C(N3086) );
and3_1 U2241 ( .Z(N7697), .A(N7531), .B(N1731), .C(N3086) );
or2_1 U2242 ( .Z(N7698), .A(N7624), .B(N7625) );
inv_1 U2243 ( .Z(N7699), .A(N7573) );
inv_1 U2244 ( .Z(N7700), .A(N7567) );
inv_1 U2245 ( .Z(N7701), .A(N7561) );
inv_1 U2246 ( .Z(N7702), .A(N7555) );
and3_1 U2247 ( .Z(N7703), .A(N1156), .B(N7631), .C(N245) );
inv_1 U2248 ( .Z(N7704), .A(N7549) );
inv_1 U2249 ( .Z(N7705), .A(N7543) );
inv_1 U2250 ( .Z(N7706), .A(N7537) );
inv_1 U2251 ( .Z(N7707), .A(N7531) );
inv_1 U2252 ( .Z(N7708), .A(N7579) );
nand2_1 U2253 ( .Z(N7709), .A(N7579), .B(N6739) );
inv_1 U2254 ( .Z(N7710), .A(N7582) );
nand2_1 U2255 ( .Z(N7711), .A(N7582), .B(N6744) );
nand2_1 U2256 ( .Z(N7712), .A(N7657), .B(N7586) );
nand2_1 U2257 ( .Z(N7715), .A(N7658), .B(N7588) );
inv_1 U2258 ( .Z(N7718), .A(N7589) );
nand2_1 U2259 ( .Z(N7719), .A(N7589), .B(N6772) );
inv_1 U2260 ( .Z(N7720), .A(N7592) );
nand2_1 U2261 ( .Z(N7721), .A(N7592), .B(N6776) );
inv_1 U2262 ( .Z(N7722), .A(N7595) );
nand2_1 U2263 ( .Z(N7723), .A(N7595), .B(N5733) );
nand2_1 U2264 ( .Z(N7724), .A(N7665), .B(N7599) );
or4_1 U2265 ( .Z(N7727), .A(N7666), .B(N7667), .C(N3617), .D(N2586) );
or4_1 U2266 ( .Z(N7728), .A(N7668), .B(N7669), .C(N3618), .D(N2587) );
or4_1 U2267 ( .Z(N7729), .A(N7670), .B(N7671), .C(N3619), .D(N2588) );
or4_1 U2268 ( .Z(N7730), .A(N7672), .B(N7673), .C(N3620), .D(N2589) );
or4_1 U2269 ( .Z(N7731), .A(N7674), .B(N7675), .C(N3628), .D(N2596) );
or4_1 U2270 ( .Z(N7732), .A(N7676), .B(N7677), .C(N3629), .D(N2597) );
or4_1 U2271 ( .Z(N7733), .A(N7678), .B(N7679), .C(N3630), .D(N2598) );
or4_1 U2272 ( .Z(N7734), .A(N7680), .B(N7681), .C(N3631), .D(N2599) );
or4_1 U2273 ( .Z(N7735), .A(N7682), .B(N7683), .C(N3638), .D(N2604) );
or4_1 U2274 ( .Z(N7736), .A(N7684), .B(N7685), .C(N3642), .D(N2606) );
or4_1 U2275 ( .Z(N7737), .A(N7686), .B(N7687), .C(N3643), .D(N2607) );
or4_1 U2276 ( .Z(N7738), .A(N7688), .B(N7689), .C(N3644), .D(N2608) );
or4_1 U2277 ( .Z(N7739), .A(N7690), .B(N7691), .C(N3645), .D(N2609) );
or4_1 U2278 ( .Z(N7740), .A(N7692), .B(N7693), .C(N3651), .D(N2615) );
or4_1 U2279 ( .Z(N7741), .A(N7694), .B(N7695), .C(N3652), .D(N2616) );
or4_1 U2280 ( .Z(N7742), .A(N7696), .B(N7697), .C(N3653), .D(N2617) );
nand2_1 U2281 ( .Z(N7743), .A(N6271), .B(N7708) );
nand2_1 U2282 ( .Z(N7744), .A(N6283), .B(N7710) );
nand2_1 U2283 ( .Z(N7749), .A(N6341), .B(N7718) );
nand2_1 U2284 ( .Z(N7750), .A(N6347), .B(N7720) );
nand2_1 U2285 ( .Z(N7751), .A(N5214), .B(N7722) );
and2_1 U2286 ( .Z(N7754), .A(N7727), .B(N2647) );
and2_1 U2287 ( .Z(N7755), .A(N7728), .B(N2647) );
and2_1 U2288 ( .Z(N7756), .A(N7729), .B(N2647) );
and2_1 U2289 ( .Z(N7757), .A(N7730), .B(N2647) );
and2_1 U2290 ( .Z(N7758), .A(N7731), .B(N2722) );
and2_1 U2291 ( .Z(N7759), .A(N7732), .B(N2722) );
and2_1 U2292 ( .Z(N7760), .A(N7733), .B(N2722) );
and2_1 U2293 ( .Z(N7761), .A(N7734), .B(N2722) );
nand2_1 U2294 ( .Z(N7762), .A(N7743), .B(N7709) );
nand2_1 U2295 ( .Z(N7765), .A(N7744), .B(N7711) );
inv_1 U2296 ( .Z(N7768), .A(N7712) );
nand2_1 U2297 ( .Z(N7769), .A(N7712), .B(N6751) );
inv_1 U2298 ( .Z(N7770), .A(N7715) );
nand2_1 U2299 ( .Z(N7771), .A(N7715), .B(N6760) );
nand2_1 U2300 ( .Z(N7772), .A(N7749), .B(N7719) );
nand2_1 U2301 ( .Z(N7775), .A(N7750), .B(N7721) );
nand2_1 U2302 ( .Z(N7778), .A(N7751), .B(N7723) );
inv_1 U2303 ( .Z(N7781), .A(N7724) );
nand2_1 U2304 ( .Z(N7782), .A(N7724), .B(N5735) );
nand2_1 U2305 ( .Z(N7787), .A(N6295), .B(N7768) );
nand2_1 U2306 ( .Z(N7788), .A(N6313), .B(N7770) );
nand2_1 U2307 ( .Z(N7795), .A(N5220), .B(N7781) );
inv_1 U2308 ( .Z(N7796), .A(N7762) );
nand2_1 U2309 ( .Z(N7797), .A(N7762), .B(N6740) );
inv_1 U2310 ( .Z(N7798), .A(N7765) );
nand2_1 U2311 ( .Z(N7799), .A(N7765), .B(N6745) );
nand2_1 U2312 ( .Z(N7800), .A(N7787), .B(N7769) );
nand2_1 U2313 ( .Z(N7803), .A(N7788), .B(N7771) );
inv_1 U2314 ( .Z(N7806), .A(N7772) );
nand2_1 U2315 ( .Z(N7807), .A(N7772), .B(N6773) );
inv_1 U2316 ( .Z(N7808), .A(N7775) );
nand2_1 U2317 ( .Z(N7809), .A(N7775), .B(N6777) );
inv_1 U2318 ( .Z(N7810), .A(N7778) );
nand2_1 U2319 ( .Z(N7811), .A(N7778), .B(N6782) );
nand2_1 U2320 ( .Z(N7812), .A(N7795), .B(N7782) );
nand2_1 U2321 ( .Z(N7815), .A(N6274), .B(N7796) );
nand2_1 U2322 ( .Z(N7816), .A(N6286), .B(N7798) );
nand2_1 U2323 ( .Z(N7821), .A(N6344), .B(N7806) );
nand2_1 U2324 ( .Z(N7822), .A(N6350), .B(N7808) );
nand2_1 U2325 ( .Z(N7823), .A(N6353), .B(N7810) );
nand2_1 U2326 ( .Z(N7826), .A(N7815), .B(N7797) );
nand2_1 U2327 ( .Z(N7829), .A(N7816), .B(N7799) );
inv_1 U2328 ( .Z(N7832), .A(N7800) );
nand2_1 U2329 ( .Z(N7833), .A(N7800), .B(N6752) );
inv_1 U2330 ( .Z(N7834), .A(N7803) );
nand2_1 U2331 ( .Z(N7835), .A(N7803), .B(N6761) );
nand2_1 U2332 ( .Z(N7836), .A(N7821), .B(N7807) );
nand2_1 U2333 ( .Z(N7839), .A(N7822), .B(N7809) );
nand2_1 U2334 ( .Z(N7842), .A(N7823), .B(N7811) );
inv_1 U2335 ( .Z(N7845), .A(N7812) );
nand2_1 U2336 ( .Z(N7846), .A(N7812), .B(N6790) );
nand2_1 U2337 ( .Z(N7851), .A(N6298), .B(N7832) );
nand2_1 U2338 ( .Z(N7852), .A(N6316), .B(N7834) );
nand2_1 U2339 ( .Z(N7859), .A(N6364), .B(N7845) );
inv_1 U2340 ( .Z(N7860), .A(N7826) );
nand2_1 U2341 ( .Z(N7861), .A(N7826), .B(N6741) );
inv_1 U2342 ( .Z(N7862), .A(N7829) );
nand2_1 U2343 ( .Z(N7863), .A(N7829), .B(N6746) );
nand2_1 U2344 ( .Z(N7864), .A(N7851), .B(N7833) );
nand2_1 U2345 ( .Z(N7867), .A(N7852), .B(N7835) );
inv_1 U2346 ( .Z(N7870), .A(N7836) );
nand2_1 U2347 ( .Z(N7871), .A(N7836), .B(N5730) );
inv_1 U2348 ( .Z(N7872), .A(N7839) );
nand2_1 U2349 ( .Z(N7873), .A(N7839), .B(N5732) );
inv_1 U2350 ( .Z(N7874), .A(N7842) );
nand2_1 U2351 ( .Z(N7875), .A(N7842), .B(N6783) );
nand2_1 U2352 ( .Z(N7876), .A(N7859), .B(N7846) );
nand2_1 U2353 ( .Z(N7879), .A(N6277), .B(N7860) );
nand2_1 U2354 ( .Z(N7880), .A(N6289), .B(N7862) );
nand2_1 U2355 ( .Z(N7885), .A(N5199), .B(N7870) );
nand2_1 U2356 ( .Z(N7886), .A(N5208), .B(N7872) );
nand2_1 U2357 ( .Z(N7887), .A(N6356), .B(N7874) );
nand2_1 U2358 ( .Z(N7890), .A(N7879), .B(N7861) );
nand2_1 U2359 ( .Z(N7893), .A(N7880), .B(N7863) );
inv_1 U2360 ( .Z(N7896), .A(N7864) );
nand2_1 U2361 ( .Z(N7897), .A(N7864), .B(N6753) );
inv_1 U2362 ( .Z(N7898), .A(N7867) );
nand2_1 U2363 ( .Z(N7899), .A(N7867), .B(N6762) );
nand2_1 U2364 ( .Z(N7900), .A(N7885), .B(N7871) );
nand2_1 U2365 ( .Z(N7903), .A(N7886), .B(N7873) );
nand2_1 U2366 ( .Z(N7906), .A(N7887), .B(N7875) );
inv_1 U2367 ( .Z(N7909), .A(N7876) );
nand2_1 U2368 ( .Z(N7910), .A(N7876), .B(N6791) );
nand2_1 U2369 ( .Z(N7917), .A(N6301), .B(N7896) );
nand2_1 U2370 ( .Z(N7918), .A(N6319), .B(N7898) );
nand2_1 U2371 ( .Z(N7923), .A(N6367), .B(N7909) );
inv_1 U2372 ( .Z(N7924), .A(N7890) );
nand2_1 U2373 ( .Z(N7925), .A(N7890), .B(N6680) );
inv_1 U2374 ( .Z(N7926), .A(N7893) );
nand2_1 U2375 ( .Z(N7927), .A(N7893), .B(N6681) );
inv_1 U2376 ( .Z(N7928), .A(N7900) );
nand2_1 U2377 ( .Z(N7929), .A(N7900), .B(N5690) );
inv_1 U2378 ( .Z(N7930), .A(N7903) );
nand2_1 U2379 ( .Z(N7931), .A(N7903), .B(N5691) );
nand2_1 U2380 ( .Z(N7932), .A(N7917), .B(N7897) );
nand2_1 U2381 ( .Z(N7935), .A(N7918), .B(N7899) );
inv_1 U2382 ( .Z(N7938), .A(N7906) );
nand2_1 U2383 ( .Z(N7939), .A(N7906), .B(N6784) );
nand2_1 U2384 ( .Z(N7940), .A(N7923), .B(N7910) );
nand2_1 U2385 ( .Z(N7943), .A(N6280), .B(N7924) );
nand2_1 U2386 ( .Z(N7944), .A(N6292), .B(N7926) );
nand2_1 U2387 ( .Z(N7945), .A(N5202), .B(N7928) );
nand2_1 U2388 ( .Z(N7946), .A(N5211), .B(N7930) );
nand2_1 U2389 ( .Z(N7951), .A(N6359), .B(N7938) );
nand2_1 U2390 ( .Z(N7954), .A(N7943), .B(N7925) );
nand2_1 U2391 ( .Z(N7957), .A(N7944), .B(N7927) );
nand2_1 U2392 ( .Z(N7960), .A(N7945), .B(N7929) );
nand2_1 U2393 ( .Z(N7963), .A(N7946), .B(N7931) );
inv_1 U2394 ( .Z(N7966), .A(N7932) );
nand2_1 U2395 ( .Z(N7967), .A(N7932), .B(N6754) );
inv_1 U2396 ( .Z(N7968), .A(N7935) );
nand2_1 U2397 ( .Z(N7969), .A(N7935), .B(N6755) );
nand2_1 U2398 ( .Z(N7970), .A(N7951), .B(N7939) );
inv_1 U2399 ( .Z(N7973), .A(N7940) );
nand2_1 U2400 ( .Z(N7974), .A(N7940), .B(N6785) );
nand2_1 U2401 ( .Z(N7984), .A(N6304), .B(N7966) );
nand2_1 U2402 ( .Z(N7985), .A(N6322), .B(N7968) );
nand2_1 U2403 ( .Z(N7987), .A(N6370), .B(N7973) );
and3_1 U2404 ( .Z(N7988), .A(N7957), .B(N6831), .C(N1157) );
and3_1 U2405 ( .Z(N7989), .A(N7954), .B(N6415), .C(N1157) );
and3_1 U2406 ( .Z(N7990), .A(N7957), .B(N7041), .C(N566) );
and3_1 U2407 ( .Z(N7991), .A(N7954), .B(N7177), .C(N566) );
inv_1 U2408 ( .Z(N7992), .A(N7970) );
nand2_1 U2409 ( .Z(N7993), .A(N7970), .B(N6448) );
and3_1 U2410 ( .Z(N7994), .A(N7963), .B(N6857), .C(N1219) );
and3_1 U2411 ( .Z(N7995), .A(N7960), .B(N6441), .C(N1219) );
and3_1 U2412 ( .Z(N7996), .A(N7963), .B(N7065), .C(N583) );
and3_1 U2413 ( .Z(N7997), .A(N7960), .B(N7182), .C(N583) );
nand2_1 U2414 ( .Z(N7998), .A(N7984), .B(N7967) );
nand2_1 U2415 ( .Z(N8001), .A(N7985), .B(N7969) );
nand2_1 U2416 ( .Z(N8004), .A(N7987), .B(N7974) );
nand2_1 U2417 ( .Z(N8009), .A(N6051), .B(N7992) );
or4_1 U2418 ( .Z(N8013), .A(N7988), .B(N7989), .C(N7990), .D(N7991) );
or4_1 U2419 ( .Z(N8017), .A(N7994), .B(N7995), .C(N7996), .D(N7997) );
inv_1 U2420 ( .Z(N8020), .A(N7998) );
nand2_1 U2421 ( .Z(N8021), .A(N7998), .B(N6682) );
inv_1 U2422 ( .Z(N8022), .A(N8001) );
nand2_1 U2423 ( .Z(N8023), .A(N8001), .B(N6683) );
nand2_1 U2424 ( .Z(N8025), .A(N8009), .B(N7993) );
inv_1 U2425 ( .Z(N8026), .A(N8004) );
nand2_1 U2426 ( .Z(N8027), .A(N8004), .B(N6449) );
nand2_1 U2427 ( .Z(N8031), .A(N6307), .B(N8020) );
nand2_1 U2428 ( .Z(N8032), .A(N6310), .B(N8022) );
inv_1 U2429 ( .Z(N8033), .A(N8013) );
nand2_1 U2430 ( .Z(N8034), .A(N6054), .B(N8026) );
and2_1 U2431 ( .Z(N8035), .A(N583), .B(N8025) );
inv_1 U2432 ( .Z(N8036), .A(N8017) );
nand2_1 U2433 ( .Z(N8037), .A(N8031), .B(N8021) );
nand2_1 U2434 ( .Z(N8038), .A(N8032), .B(N8023) );
nand2_1 U2435 ( .Z(N8039), .A(N8034), .B(N8027) );
inv_1 U2436 ( .Z(N8040), .A(N8038) );
and2_1 U2437 ( .Z(N8041), .A(N566), .B(N8037) );
inv_1 U2438 ( .Z(N8042), .A(N8039) );
and2_1 U2439 ( .Z(N8043), .A(N8040), .B(N1157) );
and2_1 U2440 ( .Z(N8044), .A(N8042), .B(N1219) );
or2_1 U2441 ( .Z(N8045), .A(N8043), .B(N8041) );
or2_1 U2442 ( .Z(N8048), .A(N8044), .B(N8035) );
nand2_1 U2443 ( .Z(N8055), .A(N8045), .B(N8033) );
inv_1 U2444 ( .Z(N8056), .A(N8045) );
nand2_1 U2445 ( .Z(N8057), .A(N8048), .B(N8036) );
inv_1 U2446 ( .Z(N8058), .A(N8048) );
nand2_1 U2447 ( .Z(N8059), .A(N8013), .B(N8056) );
nand2_1 U2448 ( .Z(N8060), .A(N8017), .B(N8058) );
nand2_1 U2449 ( .Z(N8061), .A(N8055), .B(N8059) );
nand2_1 U2450 ( .Z(N8064), .A(N8057), .B(N8060) );
and3_1 U2451 ( .Z(N8071), .A(N8064), .B(N1777), .C(N3130) );
and3_1 U2452 ( .Z(N8072), .A(N8061), .B(N1761), .C(N3108) );
inv_1 U2453 ( .Z(N8073), .A(N8061) );
inv_1 U2454 ( .Z(N8074), .A(N8064) );
or4_1 U2455 ( .Z(N8075), .A(N7526), .B(N8071), .C(N3659), .D(N2625) );
or4_1 U2456 ( .Z(N8076), .A(N7636), .B(N8072), .C(N3661), .D(N2627) );
and2_1 U2457 ( .Z(N8077), .A(N8073), .B(N1727) );
and2_1 U2458 ( .Z(N8078), .A(N8074), .B(N1727) );
or2_1 U2459 ( .Z(N8079), .A(N7530), .B(N8077) );
or2_1 U2460 ( .Z(N8082), .A(N7479), .B(N8078) );
and2_1 U2461 ( .Z(N8089), .A(N8079), .B(N3063) );
and2_1 U2462 ( .Z(N8090), .A(N8082), .B(N3063) );
and2_1 U2463 ( .Z(N8091), .A(N8079), .B(N3063) );
and2_1 U2464 ( .Z(N8092), .A(N8082), .B(N3063) );
or2_1 U2465 ( .Z(N8093), .A(N8089), .B(N3071) );
or2_1 U2466 ( .Z(N8096), .A(N8090), .B(N3072) );
or2_1 U2467 ( .Z(N8099), .A(N8091), .B(N3073) );
or2_1 U2468 ( .Z(N8102), .A(N8092), .B(N3074) );
and3_1 U2469 ( .Z(N8113), .A(N8102), .B(N2779), .C(N2790) );
and3_1 U2470 ( .Z(N8114), .A(N8099), .B(N1327), .C(N2790) );
and3_1 U2471 ( .Z(N8115), .A(N8102), .B(N2801), .C(N2812) );
and3_1 U2472 ( .Z(N8116), .A(N8099), .B(N1351), .C(N2812) );
and3_1 U2473 ( .Z(N8117), .A(N8096), .B(N2681), .C(N2692) );
and3_1 U2474 ( .Z(N8118), .A(N8093), .B(N1185), .C(N2692) );
and3_1 U2475 ( .Z(N8119), .A(N8096), .B(N2756), .C(N2767) );
and3_1 U2476 ( .Z(N8120), .A(N8093), .B(N1247), .C(N2767) );
or4_1 U2477 ( .Z(N8121), .A(N8117), .B(N8118), .C(N3662), .D(N2703) );
or4_1 U2478 ( .Z(N8122), .A(N8119), .B(N8120), .C(N3663), .D(N2778) );
or4_1 U2479 ( .Z(N8123), .A(N8113), .B(N8114), .C(N3650), .D(N2614) );
or4_1 U2480 ( .Z(N8124), .A(N8115), .B(N8116), .C(N3658), .D(N2622) );
and2_1 U2481 ( .Z(N8125), .A(N8121), .B(N2675) );
and2_1 U2482 ( .Z(N8126), .A(N8122), .B(N2750) );
inv_1 U2483 ( .Z(N8127), .A(N8125) );
inv_1 U2484 ( .Z(N8128), .A(N8126) );

endmodule
