`timescale 1ns / 1ps

module amux (
  // Mux Inputs
  input   logic [7:0] Cnt1_Out,
  input   logic [7:0] Cnt2_Out,
  // Mux Selection
  input   logic       Sel_Mux,
  // Mux Output
  output  logic [7:0] Mux_Addr
);

////////////////////////////////////////////////////////////////
///////////////////////   Module Logic   ///////////////////////
////////////////////////////////////////////////////////////////

assign Mux_Addr = (Sel_Mux == 1'b1) ? Cnt2_Out : Cnt1_Out;

////////////////////////////////////////////////////////////////
//////////////////   Instantiation Template   //////////////////
////////////////////////////////////////////////////////////////
/*
amux amux (
  .Cnt1_Out(),
  .Cnt2_Out(),
  .Sel_Mux(),
  .Mux_Addr()
);
*/
endmodule