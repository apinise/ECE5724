module mem_buffer (
  // Clk + Reset
  input   logic         Clk,
  input   logic         Rst,
  // Read + Write Ctrl
  input   logic         Read,
  input   logic         Write,
  // Read + Write Ports
  input   logic [7:0]   Address,
  input   logic [15:0]  Write_Data,
  output  logic [15:0]  Read_Data
);

////////////////////////////////////////////////////////////////
////////////////////////   Parameters   ////////////////////////
////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////
///////////////////////   Internal Net   ///////////////////////
////////////////////////////////////////////////////////////////

logic [15:0]  data_mem  [255:0];

////////////////////////////////////////////////////////////////
//////////////////////   Instantiations   //////////////////////
////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////
///////////////////////   Module Logic   ///////////////////////
////////////////////////////////////////////////////////////////

initial begin
  $readmemb("./data.txt", data_mem);
end

// Write Port
always_ff @(posedge Clk) begin
  if (Rst) begin
    $readmemb("./data.txt", data_mem);
  end
  else begin
    if (Write) begin
      data_mem[Address] <= Write_Data;
    end
  end
end

// Read Port
always_ff @(posedge Clk) begin
  if (Rst) begin
    Read_Data <= '0;
  end
  else begin
    if (Read) begin
      Read_Data <= data_mem[Address];
    end
    else begin
      Read_Data <= 'z;
    end
  end
end

////////////////////////////////////////////////////////////////
//////////////////   Instantiation Template   //////////////////
////////////////////////////////////////////////////////////////

endmodule