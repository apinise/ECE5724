`timescale 1ns / 1ps

module data_mux (
  // Mux Inputs
  input   logic [15:0]  Min_Reg,
  input   logic [15:0]  Temp_Reg,
  // Mux Selection
  input   logic         Sel_DMux,
  // Mux Output To Mem Buffer
  output  logic [15:0]  Write_Data
);

////////////////////////////////////////////////////////////////
///////////////////////   Module Logic   ///////////////////////
////////////////////////////////////////////////////////////////

assign Write_Data = Sel_DMux ? Temp_Reg : Min_Reg;

////////////////////////////////////////////////////////////////
//////////////////   Instantiation Template   //////////////////
////////////////////////////////////////////////////////////////
/*
data_mux data_mux (
  .Min_Reg(),
  .Temp_Reg(),
  .Sel_DMux(),
  .Write_Data()
);
*/
endmodule