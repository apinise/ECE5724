
//Verilog file of module SSC


`timescale 1 ns / 1ns

module SSC_net(clk,
rst,
start,
read_reg,
write_reg,
readdata,
writedata,
addr,
done,
Si,
So,
NbarT);
	input clk;
	input rst;
	input start;
  input [0:15]readdata;
  input NbarT, Si;

  output So;
  output [0:15]writedata;
  output [0:7]addr;
	output read_reg;
	output write_reg;
	output done;

wire
SSC_wire_1,
SSC_wire_2,
SSC_wire_3,
SSC_wire_4,
SSC_wire_5,
SSC_wire_6,
SSC_wire_7,
SSC_wire_8,
SSC_wire_9,
SSC_wire_10,
SSC_wire_11,
SSC_wire_12,
SSC_wire_13,
SSC_wire_14,
SSC_wire_15,
SSC_wire_16,
SSC_wire_17,
SSC_wire_18,
SSC_wire_19,
SSC_wire_20,
SSC_wire_21,
SSC_wire_22,
SSC_wire_23,
SSC_wire_24,
SSC_wire_25,
SSC_wire_26,
SSC_wire_27,
SSC_wire_28,
SSC_wire_29,
SSC_wire_30,
SSC_wire_31,
SSC_wire_32,
SSC_wire_33,
SSC_wire_34,
SSC_wire_35,
SSC_wire_36,
SSC_wire_37,
SSC_wire_38,
SSC_wire_39,
SSC_wire_40,
SSC_wire_41,
SSC_wire_42,
SSC_wire_43,
SSC_wire_44,
SSC_wire_45,
SSC_wire_46,
SSC_wire_47,
SSC_wire_48,
SSC_wire_49,
SSC_wire_50,
SSC_wire_51,
SSC_wire_52,
SSC_wire_53,
SSC_wire_54,
SSC_wire_55,
SSC_wire_56,
SSC_wire_57,
SSC_wire_58,
SSC_wire_59,
SSC_wire_60,
SSC_wire_61,
SSC_wire_62,
SSC_wire_63,
SSC_wire_64,
SSC_wire_65,
SSC_wire_66,
SSC_wire_67,
SSC_wire_68,
SSC_wire_69,
SSC_wire_70,
SSC_wire_71,
SSC_wire_72,
SSC_wire_73,
SSC_wire_74,
SSC_wire_75,
SSC_wire_76,
SSC_wire_77,
SSC_wire_78,
SSC_wire_79,
SSC_wire_80,
SSC_wire_81,
SSC_wire_82,
SSC_wire_83,
SSC_wire_84,
SSC_wire_85,
SSC_wire_86,
SSC_wire_87,
SSC_wire_88,
SSC_wire_89,
SSC_wire_90,
SSC_wire_91,
SSC_wire_92,
SSC_wire_93,
SSC_wire_94,
SSC_wire_95,
SSC_wire_96,
SSC_wire_97,
SSC_wire_98,
SSC_wire_99,
SSC_wire_100,
SSC_wire_101,
SSC_wire_102,
SSC_wire_103,
SSC_wire_104,
SSC_wire_105,
SSC_wire_106,
SSC_wire_107,
SSC_wire_108,
SSC_wire_109,
SSC_wire_110,
SSC_wire_111,
SSC_wire_112,
SSC_wire_113,
SSC_wire_114,
SSC_wire_115,
SSC_wire_116,
SSC_wire_117,
SSC_wire_118,
SSC_wire_119,
SSC_wire_120,
SSC_wire_121,
SSC_wire_122,
SSC_wire_123,
SSC_wire_124,
SSC_wire_125,
SSC_wire_126,
SSC_wire_127,
SSC_wire_128,
SSC_wire_129,
SSC_wire_130,
SSC_wire_131,
SSC_wire_132,
SSC_wire_133,
SSC_wire_134,
SSC_wire_135,
SSC_wire_136,
SSC_wire_137,
SSC_wire_138,
SSC_wire_139,
SSC_wire_140,
SSC_wire_141,
SSC_wire_142,
SSC_wire_143,
SSC_wire_144,
SSC_wire_145,
SSC_wire_146,
SSC_wire_147,
SSC_wire_148,
SSC_wire_149,
SSC_wire_150,
SSC_wire_151,
SSC_wire_152,
SSC_wire_153,
SSC_wire_154,
SSC_wire_155,
SSC_wire_156,
SSC_wire_157,
SSC_wire_158,
SSC_wire_159,
SSC_wire_160,
SSC_wire_161,
SSC_wire_162,
SSC_wire_163,
SSC_wire_164,
SSC_wire_165,
SSC_wire_166,
SSC_wire_167,
SSC_wire_168,
SSC_wire_169,
SSC_wire_170,
SSC_wire_171,
SSC_wire_172,
SSC_wire_173,
SSC_wire_174,
SSC_wire_175,
SSC_wire_176,
SSC_wire_177,
SSC_wire_178,
SSC_wire_179,
SSC_wire_180,
SSC_wire_181,
SSC_wire_182,
SSC_wire_183,
SSC_wire_184,
SSC_wire_185,
SSC_wire_186,
SSC_wire_187,
SSC_wire_188,
SSC_wire_189,
SSC_wire_190,
SSC_wire_191,
SSC_wire_192,
SSC_wire_193,
SSC_wire_194,
SSC_wire_195,
SSC_wire_196,
SSC_wire_197,
SSC_wire_198,
SSC_wire_199,
SSC_wire_200,
SSC_wire_201,
SSC_wire_202,
SSC_wire_203,
SSC_wire_204,
SSC_wire_205,
SSC_wire_206,
SSC_wire_207,
SSC_wire_208,
SSC_wire_209,
SSC_wire_210,
SSC_wire_211,
SSC_wire_212,
SSC_wire_213,
SSC_wire_214,
SSC_wire_215,
SSC_wire_216,
SSC_wire_217,
SSC_wire_218,
SSC_wire_219,
SSC_wire_220,
SSC_wire_221,
SSC_wire_222,
SSC_wire_223,
SSC_wire_224,
SSC_wire_225,
SSC_wire_226,
SSC_wire_227,
SSC_wire_228,
SSC_wire_229,
SSC_wire_230,
SSC_wire_231,
SSC_wire_232,
SSC_wire_233,
SSC_wire_234,
SSC_wire_235,
SSC_wire_236,
SSC_wire_237,
SSC_wire_238,
SSC_wire_239,
SSC_wire_240,
SSC_wire_241,
SSC_wire_242,
SSC_wire_243,
SSC_wire_244,
SSC_wire_245,
SSC_wire_246,
SSC_wire_247,
SSC_wire_248,
SSC_wire_249,
SSC_wire_250,
SSC_wire_251,
SSC_wire_252,
SSC_wire_253,
SSC_wire_254,
SSC_wire_255,
SSC_wire_256,
SSC_wire_257,
SSC_wire_258,
SSC_wire_259,
SSC_wire_260,
SSC_wire_261,
SSC_wire_262,
SSC_wire_263,
SSC_wire_264,
SSC_wire_265,
SSC_wire_266,
SSC_wire_267,
SSC_wire_268,
SSC_wire_269,
SSC_wire_270,
SSC_wire_271,
SSC_wire_272,
SSC_wire_273,
SSC_wire_274,
SSC_wire_275,
SSC_wire_276,
SSC_wire_277,
SSC_wire_278,
SSC_wire_279,
SSC_wire_280,
SSC_wire_281,
SSC_wire_282,
SSC_wire_283,
SSC_wire_284,
SSC_wire_285,
SSC_wire_286,
SSC_wire_287,
SSC_wire_288,
SSC_wire_289,
SSC_wire_290,
SSC_wire_291,
SSC_wire_292,
SSC_wire_293,
SSC_wire_294,
SSC_wire_295,
SSC_wire_296,
SSC_wire_297,
SSC_wire_298,
SSC_wire_299,
SSC_wire_300,
SSC_wire_301,
SSC_wire_302,
SSC_wire_303,
SSC_wire_304,
SSC_wire_305,
SSC_wire_306,
SSC_wire_307,
SSC_wire_308,
SSC_wire_309,
SSC_wire_310,
SSC_wire_311,
SSC_wire_312,
SSC_wire_313,
SSC_wire_314,
SSC_wire_315,
SSC_wire_316,
SSC_wire_317,
SSC_wire_318,
SSC_wire_319,
SSC_wire_320,
SSC_wire_321,
SSC_wire_322,
SSC_wire_323,
SSC_wire_324,
SSC_wire_325,
SSC_wire_326,
SSC_wire_327,
SSC_wire_328,
SSC_wire_329,
SSC_wire_330,
SSC_wire_331,
SSC_wire_332,
SSC_wire_333,
SSC_wire_334,
SSC_wire_335,
SSC_wire_336,
SSC_wire_337,
SSC_wire_338,
SSC_wire_339,
SSC_wire_340,
SSC_wire_341,
SSC_wire_342,
SSC_wire_343,
SSC_wire_344,
SSC_wire_345,
SSC_wire_346,
SSC_wire_347,
SSC_wire_348,
SSC_wire_349,
SSC_wire_350,
SSC_wire_351,
SSC_wire_352,
SSC_wire_353,
SSC_wire_354,
SSC_wire_355,
SSC_wire_356,
SSC_wire_357,
SSC_wire_358,
SSC_wire_359,
SSC_wire_360,
SSC_wire_361,
SSC_wire_362,
SSC_wire_363,
SSC_wire_364,
SSC_wire_365,
SSC_wire_366,
SSC_wire_367,
SSC_wire_368,
SSC_wire_369,
SSC_wire_370,
SSC_wire_371,
SSC_wire_372,
SSC_wire_373,
SSC_wire_374,
SSC_wire_375,
SSC_wire_376,
SSC_wire_377,
SSC_wire_378,
SSC_wire_379,
SSC_wire_380,
SSC_wire_381,
SSC_wire_382,
SSC_wire_383,
SSC_wire_384,
SSC_wire_385,
SSC_wire_386,
SSC_wire_387,
SSC_wire_388,
SSC_wire_389,
SSC_wire_390,
SSC_wire_391,
SSC_wire_392,
SSC_wire_393,
SSC_wire_394,
SSC_wire_395,
SSC_wire_396,
SSC_wire_397,
SSC_wire_398,
SSC_wire_399,
SSC_wire_400,
SSC_wire_401,
SSC_wire_402,
SSC_wire_403,
SSC_wire_404,
SSC_wire_405,
SSC_wire_406,
SSC_wire_407,
SSC_wire_408,
SSC_wire_409,
SSC_wire_410,
SSC_wire_411,
SSC_wire_412,
SSC_wire_413,
SSC_wire_414,
SSC_wire_415,
SSC_wire_416,
SSC_wire_417,
SSC_wire_418,
SSC_wire_419,
SSC_wire_420,
SSC_wire_421,
SSC_wire_422,
SSC_wire_423,
SSC_wire_424,
SSC_wire_425,
SSC_wire_426,
SSC_wire_427,
SSC_wire_428,
SSC_wire_429,
SSC_wire_430,
SSC_wire_431,
SSC_wire_432,
SSC_wire_433,
SSC_wire_434,
SSC_wire_435,
SSC_wire_436,
SSC_wire_437,
SSC_wire_438,
SSC_wire_439,
SSC_wire_440,
SSC_wire_441,
SSC_wire_442,
SSC_wire_443,
SSC_wire_444,
SSC_wire_445,
SSC_wire_446,
SSC_wire_447,
SSC_wire_448,
SSC_wire_449,
SSC_wire_450,
SSC_wire_451,
SSC_wire_452,
SSC_wire_453,
SSC_wire_454,
SSC_wire_455,
SSC_wire_456,
SSC_wire_457,
SSC_wire_458,
SSC_wire_459,
SSC_wire_460,
SSC_wire_461,
SSC_wire_462,
SSC_wire_463,
SSC_wire_464,
SSC_wire_465,
SSC_wire_466,
SSC_wire_467,
SSC_wire_468,
SSC_wire_469,
SSC_wire_470,
SSC_wire_471,
SSC_wire_472,
SSC_wire_473,
SSC_wire_474,
SSC_wire_475,
SSC_wire_476,
SSC_wire_477,
SSC_wire_478,
SSC_wire_479,
SSC_wire_480,
SSC_wire_481,
SSC_wire_482,
SSC_wire_483,
SSC_wire_484,
SSC_wire_485,
SSC_wire_486,
SSC_wire_487,
SSC_wire_488,
SSC_wire_489,
SSC_wire_490,
SSC_wire_491,
SSC_wire_492,
SSC_wire_493,
SSC_wire_494,
SSC_wire_495,
SSC_wire_496,
SSC_wire_497,
SSC_wire_498,
SSC_wire_499,
SSC_wire_500,
SSC_wire_501,
SSC_wire_502,
SSC_wire_503,
SSC_wire_504,
SSC_wire_505,
SSC_wire_506,
SSC_wire_507,
SSC_wire_508,
SSC_wire_509,
SSC_wire_510,
SSC_wire_511,
SSC_wire_73_0,
SSC_wire_73_1,
SSC_wire_73_2,
SSC_wire_73_3,
SSC_wire_73_4,
SSC_wire_73_5,
SSC_wire_71_0,
SSC_wire_71_1,
SSC_wire_71_2,
SSC_wire_71_3,
SSC_wire_71_4,
SSC_wire_69_0,
SSC_wire_69_1,
SSC_wire_69_2,
SSC_wire_69_3,
SSC_wire_67_0,
SSC_wire_67_1,
SSC_wire_67_2,
SSC_wire_67_3,
SSC_wire_65_0,
SSC_wire_65_1,
SSC_wire_65_2,
SSC_wire_65_3,
SSC_wire_63_0,
SSC_wire_63_1,
SSC_wire_63_2,
SSC_wire_63_3,
SSC_wire_91_0,
SSC_wire_91_1,
SSC_wire_91_2,
SSC_wire_89_0,
SSC_wire_89_1,
SSC_wire_89_2,
SSC_wire_89_3,
SSC_wire_89_4,
SSC_wire_87_0,
SSC_wire_87_1,
SSC_wire_87_2,
SSC_wire_87_3,
SSC_wire_85_0,
SSC_wire_85_1,
SSC_wire_85_2,
SSC_wire_85_3,
SSC_wire_83_0,
SSC_wire_83_1,
SSC_wire_83_2,
SSC_wire_81_0,
SSC_wire_81_1,
SSC_wire_81_2,
SSC_wire_81_3,
SSC_wire_79_0,
SSC_wire_79_1,
SSC_wire_79_2,
SSC_wire_77_0,
SSC_wire_77_1,
SSC_wire_77_2,
SSC_wire_75_0,
SSC_wire_75_1,
SSC_wire_75_2,
SSC_wire_60_0,
SSC_wire_60_1,
SSC_wire_19_0,
SSC_wire_19_1,
SSC_wire_19_2,
SSC_wire_19_3,
SSC_wire_19_4,
SSC_wire_19_5,
SSC_wire_22_0,
SSC_wire_22_1,
SSC_wire_22_2,
SSC_wire_22_3,
SSC_wire_22_4,
SSC_wire_24_0,
SSC_wire_24_1,
SSC_wire_24_2,
SSC_wire_24_3,
SSC_wire_24_4,
SSC_wire_26_0,
SSC_wire_26_1,
SSC_wire_26_2,
SSC_wire_26_3,
SSC_wire_26_4,
SSC_wire_28_0,
SSC_wire_28_1,
SSC_wire_28_2,
SSC_wire_28_3,
SSC_wire_28_4,
SSC_wire_30_0,
SSC_wire_30_1,
SSC_wire_30_2,
SSC_wire_30_3,
SSC_wire_30_4,
SSC_wire_32_0,
SSC_wire_32_1,
SSC_wire_32_2,
SSC_wire_32_3,
SSC_wire_32_4,
SSC_wire_34_0,
SSC_wire_34_1,
SSC_wire_34_2,
SSC_wire_34_3,
SSC_wire_423_0,
SSC_wire_423_1,
SSC_wire_412_0,
SSC_wire_412_1,
SSC_wire_410_0,
SSC_wire_410_1,
SSC_wire_408_0,
SSC_wire_408_1,
SSC_wire_406_0,
SSC_wire_406_1,
SSC_wire_404_0,
SSC_wire_404_1,
SSC_wire_2_0,
SSC_wire_2_1,
SSC_wire_2_2,
SSC_wire_2_3,
SSC_wire_2_4,
SSC_wire_2_5,
SSC_wire_2_6,
SSC_wire_2_7,
SSC_wire_2_8,
SSC_wire_5_0,
SSC_wire_5_1,
SSC_wire_5_2,
SSC_wire_5_3,
SSC_wire_5_4,
SSC_wire_5_5,
SSC_wire_5_6,
SSC_wire_7_0,
SSC_wire_7_1,
SSC_wire_7_2,
SSC_wire_7_3,
SSC_wire_7_4,
SSC_wire_7_5,
SSC_wire_7_6,
SSC_wire_9_0,
SSC_wire_9_1,
SSC_wire_9_2,
SSC_wire_9_3,
SSC_wire_9_4,
SSC_wire_9_5,
SSC_wire_9_6,
SSC_wire_11_0,
SSC_wire_11_1,
SSC_wire_11_2,
SSC_wire_11_3,
SSC_wire_11_4,
SSC_wire_11_5,
SSC_wire_11_6,
SSC_wire_13_0,
SSC_wire_13_1,
SSC_wire_13_2,
SSC_wire_13_3,
SSC_wire_13_4,
SSC_wire_13_5,
SSC_wire_13_6,
SSC_wire_15_0,
SSC_wire_15_1,
SSC_wire_15_2,
SSC_wire_15_3,
SSC_wire_15_4,
SSC_wire_15_5,
SSC_wire_15_6,
SSC_wire_17_0,
SSC_wire_17_1,
SSC_wire_17_2,
SSC_wire_17_3,
SSC_wire_17_4,
SSC_wire_470_0,
SSC_wire_470_1,
SSC_wire_467_0,
SSC_wire_467_1,
SSC_wire_465_0,
SSC_wire_465_1,
SSC_wire_463_0,
SSC_wire_463_1,
SSC_wire_461_0,
SSC_wire_461_1,
SSC_wire_459_0,
SSC_wire_459_1,
SSC_wire_472_0,
SSC_wire_472_1,
SSC_wire_471_0,
SSC_wire_471_1,
SSC_wire_473_0,
SSC_wire_473_1,
SSC_wire_474_0,
SSC_wire_474_1,
SSC_wire_475_0,
SSC_wire_475_1,
SSC_wire_478_0,
SSC_wire_478_1,
SSC_wire_94_0,
SSC_wire_94_1,
SSC_wire_94_2,
SSC_wire_94_3,
SSC_wire_94_4,
SSC_wire_94_5,
SSC_wire_94_6,
SSC_wire_94_7,
SSC_wire_94_8,
SSC_wire_94_9,
SSC_wire_94_10,
SSC_wire_94_11,
SSC_wire_94_12,
SSC_wire_94_13,
SSC_wire_94_14,
SSC_wire_94_15,
SSC_wire_94_16,
SSC_wire_94_17,
SSC_wire_94_18,
SSC_wire_94_19,
SSC_wire_94_20,
SSC_wire_94_21,
SSC_wire_94_22,
SSC_wire_94_23,
SSC_wire_94_24,
SSC_wire_94_25,
SSC_wire_94_26,
SSC_wire_61_0,
SSC_wire_61_1,
SSC_wire_61_2,
SSC_wire_61_3,
SSC_wire_61_4,
SSC_wire_61_5,
SSC_wire_61_6,
SSC_wire_61_7,
SSC_wire_61_8,
SSC_wire_61_9,
SSC_wire_61_10,
SSC_wire_61_11,
SSC_wire_61_12,
SSC_wire_61_13,
SSC_wire_61_14,
SSC_wire_61_15,
SSC_wire_61_16,
SSC_wire_61_17,
SSC_wire_61_18,
SSC_wire_61_19,
SSC_wire_61_20,
SSC_wire_61_21,
SSC_wire_61_22,
SSC_wire_61_23,
SSC_wire_61_24,
SSC_wire_61_25,
SSC_wire_61_26,
SSC_wire_61_27,
SSC_wire_61_28,
SSC_wire_61_29,
SSC_wire_61_30,
SSC_wire_61_31,
SSC_wire_61_32,
SSC_wire_61_33,
SSC_wire_61_34,
SSC_wire_398_0,
SSC_wire_398_1,
SSC_wire_398_2,
SSC_wire_20_0,
SSC_wire_20_1,
SSC_wire_20_2,
SSC_wire_20_3,
SSC_wire_20_4,
SSC_wire_20_5,
SSC_wire_20_6,
SSC_wire_20_7,
SSC_wire_20_8,
SSC_wire_20_9,
SSC_wire_20_10,
SSC_wire_20_11,
SSC_wire_20_12,
SSC_wire_20_13,
SSC_wire_20_14,
SSC_wire_20_15,
SSC_wire_20_16,
SSC_wire_20_17,
SSC_wire_20_18,
SSC_wire_20_19,
SSC_wire_20_20,
SSC_wire_20_21,
SSC_wire_20_22,
SSC_wire_20_23,
SSC_wire_20_24,
SSC_wire_20_25,
SSC_wire_20_26,
SSC_wire_20_27,
SSC_wire_3_0,
SSC_wire_3_1,
SSC_wire_3_2,
SSC_wire_3_3,
SSC_wire_3_4,
SSC_wire_3_5,
SSC_wire_3_6,
SSC_wire_3_7,
SSC_wire_3_8,
SSC_wire_3_9,
SSC_wire_3_10,
SSC_wire_3_11,
SSC_wire_3_12,
SSC_wire_3_13,
SSC_wire_3_14,
SSC_wire_3_15,
SSC_wire_3_16,
SSC_wire_3_17,
SSC_wire_3_18,
SSC_wire_3_19,
SSC_wire_3_20,
SSC_wire_3_21,
SSC_wire_3_22,
SSC_wire_3_23,
SSC_wire_3_24,
SSC_wire_3_25,
SSC_wire_3_26,
SSC_wire_3_27,
SSC_wire_3_28,
SSC_wire_3_29,
SSC_wire_3_30,
SSC_wire_3_31,
SSC_wire_3_32,
SSC_wire_3_33,
SSC_wire_3_34,
SSC_wire_3_35,
SSC_wire_3_36,
SSC_wire_3_37,
SSC_wire_485_0,
SSC_wire_485_1,
SSC_wire_487_0,
SSC_wire_487_1,
SSC_wire_174_0,
SSC_wire_174_1,
SSC_wire_174_2,
SSC_wire_174_3,
SSC_wire_174_4,
SSC_wire_174_5,
SSC_wire_174_6,
SSC_wire_174_7,
SSC_wire_174_8,
SSC_wire_174_9,
SSC_wire_174_10,
SSC_wire_174_11,
SSC_wire_174_12,
SSC_wire_174_13,
SSC_wire_174_14,
SSC_wire_174_15,
SSC_wire_294_0,
SSC_wire_294_1,
SSC_wire_294_2,
SSC_wire_324_0,
SSC_wire_324_1,
SSC_wire_324_2,
SSC_wire_322_0,
SSC_wire_322_1,
SSC_wire_322_2,
SSC_wire_331_0,
SSC_wire_331_1,
SSC_wire_331_2,
SSC_wire_329_0,
SSC_wire_329_1,
SSC_wire_329_2,
SSC_wire_329_3,
SSC_wire_333_0,
SSC_wire_333_1,
SSC_wire_333_2,
SSC_wire_333_3,
SSC_wire_333_4,
SSC_wire_273_0,
SSC_wire_273_1,
SSC_wire_268_0,
SSC_wire_268_1,
SSC_wire_312_0,
SSC_wire_312_1,
SSC_wire_265_0,
SSC_wire_265_1,
SSC_wire_265_2,
SSC_wire_310_0,
SSC_wire_310_1,
SSC_wire_311_0,
SSC_wire_311_1,
SSC_wire_311_2,
SSC_wire_318_0,
SSC_wire_318_1,
SSC_wire_318_2,
SSC_wire_316_0,
SSC_wire_316_1,
SSC_wire_316_2,
SSC_wire_316_3,
SSC_wire_307_0,
SSC_wire_307_1,
SSC_wire_399_0,
SSC_wire_399_1,
SSC_wire_399_2,
SSC_wire_399_3,
SSC_wire_399_4,
SSC_wire_399_5,
SSC_wire_399_6,
SSC_wire_399_7,
SSC_wire_504_0,
SSC_wire_504_1,
SSC_wire_504_2,
clk_net_0,
rst_net_0,
start_net_0,
read_reg_net_0,
write_reg_net_0,
done_net_0;

pin #(19) pin_0 ({clk, rst, start, readdata[0], readdata[1], readdata[2], readdata[3], readdata[4], readdata[5], readdata[6], readdata[7], readdata[8], readdata[9], readdata[10], readdata[11], readdata[12], readdata[13], readdata[14], readdata[15]}, {clk_net_0, rst_net_0, start_net_0, readdata_0, readdata_1, readdata_2, readdata_3, readdata_4, readdata_5, readdata_6, readdata_7, readdata_8, readdata_9, readdata_10, readdata_11, readdata_12, readdata_13, readdata_14, readdata_15});

pout #(27) pout_0 ({writedata_0, writedata_1, writedata_2, writedata_3, writedata_4, writedata_5, writedata_6, writedata_7, writedata_8, writedata_9, writedata_10, writedata_11, writedata_12, writedata_13, writedata_14, writedata_15, addr_0, addr_1, addr_2, addr_3, addr_4, addr_5, addr_6, addr_7, read_reg_net_0, write_reg_net_0, done_net_0}, {writedata[0], writedata[1], writedata[2], writedata[3], writedata[4], writedata[5], writedata[6], writedata[7], writedata[8], writedata[9], writedata[10], writedata[11], writedata[12], writedata[13], writedata[14], writedata[15], addr[0], addr[1], addr[2], addr[3], addr[4], addr[5], addr[6], addr[7], read_reg, write_reg, done});

fanout_n #(6, 0, 0) FANOUT_1 (SSC_wire_73, {SSC_wire_73_0, SSC_wire_73_1, SSC_wire_73_2, SSC_wire_73_3, SSC_wire_73_4, SSC_wire_73_5});
fanout_n #(5, 0, 0) FANOUT_2 (SSC_wire_71, {SSC_wire_71_0, SSC_wire_71_1, SSC_wire_71_2, SSC_wire_71_3, SSC_wire_71_4});
fanout_n #(4, 0, 0) FANOUT_3 (SSC_wire_69, {SSC_wire_69_0, SSC_wire_69_1, SSC_wire_69_2, SSC_wire_69_3});
fanout_n #(4, 0, 0) FANOUT_4 (SSC_wire_67, {SSC_wire_67_0, SSC_wire_67_1, SSC_wire_67_2, SSC_wire_67_3});
fanout_n #(4, 0, 0) FANOUT_5 (SSC_wire_65, {SSC_wire_65_0, SSC_wire_65_1, SSC_wire_65_2, SSC_wire_65_3});
fanout_n #(4, 0, 0) FANOUT_6 (SSC_wire_63, {SSC_wire_63_0, SSC_wire_63_1, SSC_wire_63_2, SSC_wire_63_3});
fanout_n #(3, 0, 0) FANOUT_7 (SSC_wire_91, {SSC_wire_91_0, SSC_wire_91_1, SSC_wire_91_2});
fanout_n #(5, 0, 0) FANOUT_8 (SSC_wire_89, {SSC_wire_89_0, SSC_wire_89_1, SSC_wire_89_2, SSC_wire_89_3, SSC_wire_89_4});
fanout_n #(4, 0, 0) FANOUT_9 (SSC_wire_87, {SSC_wire_87_0, SSC_wire_87_1, SSC_wire_87_2, SSC_wire_87_3});
fanout_n #(4, 0, 0) FANOUT_10 (SSC_wire_85, {SSC_wire_85_0, SSC_wire_85_1, SSC_wire_85_2, SSC_wire_85_3});
fanout_n #(3, 0, 0) FANOUT_11 (SSC_wire_83, {SSC_wire_83_0, SSC_wire_83_1, SSC_wire_83_2});
fanout_n #(4, 0, 0) FANOUT_12 (SSC_wire_81, {SSC_wire_81_0, SSC_wire_81_1, SSC_wire_81_2, SSC_wire_81_3});
fanout_n #(3, 0, 0) FANOUT_13 (SSC_wire_79, {SSC_wire_79_0, SSC_wire_79_1, SSC_wire_79_2});
fanout_n #(3, 0, 0) FANOUT_14 (SSC_wire_77, {SSC_wire_77_0, SSC_wire_77_1, SSC_wire_77_2});
fanout_n #(3, 0, 0) FANOUT_15 (SSC_wire_75, {SSC_wire_75_0, SSC_wire_75_1, SSC_wire_75_2});
fanout_n #(2, 0, 0) FANOUT_16 (SSC_wire_60, {SSC_wire_60_0, SSC_wire_60_1});
fanout_n #(6, 0, 0) FANOUT_17 (SSC_wire_19, {SSC_wire_19_0, SSC_wire_19_1, SSC_wire_19_2, SSC_wire_19_3, SSC_wire_19_4, SSC_wire_19_5});
fanout_n #(5, 0, 0) FANOUT_18 (SSC_wire_22, {SSC_wire_22_0, SSC_wire_22_1, SSC_wire_22_2, SSC_wire_22_3, SSC_wire_22_4});
fanout_n #(5, 0, 0) FANOUT_19 (SSC_wire_24, {SSC_wire_24_0, SSC_wire_24_1, SSC_wire_24_2, SSC_wire_24_3, SSC_wire_24_4});
fanout_n #(5, 0, 0) FANOUT_20 (SSC_wire_26, {SSC_wire_26_0, SSC_wire_26_1, SSC_wire_26_2, SSC_wire_26_3, SSC_wire_26_4});
fanout_n #(5, 0, 0) FANOUT_21 (SSC_wire_28, {SSC_wire_28_0, SSC_wire_28_1, SSC_wire_28_2, SSC_wire_28_3, SSC_wire_28_4});
fanout_n #(5, 0, 0) FANOUT_22 (SSC_wire_30, {SSC_wire_30_0, SSC_wire_30_1, SSC_wire_30_2, SSC_wire_30_3, SSC_wire_30_4});
fanout_n #(5, 0, 0) FANOUT_23 (SSC_wire_32, {SSC_wire_32_0, SSC_wire_32_1, SSC_wire_32_2, SSC_wire_32_3, SSC_wire_32_4});
fanout_n #(4, 0, 0) FANOUT_24 (SSC_wire_34, {SSC_wire_34_0, SSC_wire_34_1, SSC_wire_34_2, SSC_wire_34_3});
fanout_n #(2, 0, 0) FANOUT_25 (SSC_wire_423, {SSC_wire_423_0, SSC_wire_423_1});
fanout_n #(2, 0, 0) FANOUT_26 (SSC_wire_412, {SSC_wire_412_0, SSC_wire_412_1});
fanout_n #(2, 0, 0) FANOUT_27 (SSC_wire_410, {SSC_wire_410_0, SSC_wire_410_1});
fanout_n #(2, 0, 0) FANOUT_28 (SSC_wire_408, {SSC_wire_408_0, SSC_wire_408_1});
fanout_n #(2, 0, 0) FANOUT_29 (SSC_wire_406, {SSC_wire_406_0, SSC_wire_406_1});
fanout_n #(2, 0, 0) FANOUT_30 (SSC_wire_404, {SSC_wire_404_0, SSC_wire_404_1});
fanout_n #(9, 0, 0) FANOUT_31 (SSC_wire_2, {SSC_wire_2_0, SSC_wire_2_1, SSC_wire_2_2, SSC_wire_2_3, SSC_wire_2_4, SSC_wire_2_5, SSC_wire_2_6, SSC_wire_2_7, SSC_wire_2_8});
fanout_n #(7, 0, 0) FANOUT_32 (SSC_wire_5, {SSC_wire_5_0, SSC_wire_5_1, SSC_wire_5_2, SSC_wire_5_3, SSC_wire_5_4, SSC_wire_5_5, SSC_wire_5_6});
fanout_n #(7, 0, 0) FANOUT_33 (SSC_wire_7, {SSC_wire_7_0, SSC_wire_7_1, SSC_wire_7_2, SSC_wire_7_3, SSC_wire_7_4, SSC_wire_7_5, SSC_wire_7_6});
fanout_n #(7, 0, 0) FANOUT_34 (SSC_wire_9, {SSC_wire_9_0, SSC_wire_9_1, SSC_wire_9_2, SSC_wire_9_3, SSC_wire_9_4, SSC_wire_9_5, SSC_wire_9_6});
fanout_n #(7, 0, 0) FANOUT_35 (SSC_wire_11, {SSC_wire_11_0, SSC_wire_11_1, SSC_wire_11_2, SSC_wire_11_3, SSC_wire_11_4, SSC_wire_11_5, SSC_wire_11_6});
fanout_n #(7, 0, 0) FANOUT_36 (SSC_wire_13, {SSC_wire_13_0, SSC_wire_13_1, SSC_wire_13_2, SSC_wire_13_3, SSC_wire_13_4, SSC_wire_13_5, SSC_wire_13_6});
fanout_n #(7, 0, 0) FANOUT_37 (SSC_wire_15, {SSC_wire_15_0, SSC_wire_15_1, SSC_wire_15_2, SSC_wire_15_3, SSC_wire_15_4, SSC_wire_15_5, SSC_wire_15_6});
fanout_n #(5, 0, 0) FANOUT_38 (SSC_wire_17, {SSC_wire_17_0, SSC_wire_17_1, SSC_wire_17_2, SSC_wire_17_3, SSC_wire_17_4});
fanout_n #(2, 0, 0) FANOUT_39 (SSC_wire_470, {SSC_wire_470_0, SSC_wire_470_1});
fanout_n #(2, 0, 0) FANOUT_40 (SSC_wire_467, {SSC_wire_467_0, SSC_wire_467_1});
fanout_n #(2, 0, 0) FANOUT_41 (SSC_wire_465, {SSC_wire_465_0, SSC_wire_465_1});
fanout_n #(2, 0, 0) FANOUT_42 (SSC_wire_463, {SSC_wire_463_0, SSC_wire_463_1});
fanout_n #(2, 0, 0) FANOUT_43 (SSC_wire_461, {SSC_wire_461_0, SSC_wire_461_1});
fanout_n #(2, 0, 0) FANOUT_44 (SSC_wire_459, {SSC_wire_459_0, SSC_wire_459_1});
fanout_n #(2, 0, 0) FANOUT_45 (SSC_wire_472, {SSC_wire_472_0, SSC_wire_472_1});
fanout_n #(2, 0, 0) FANOUT_46 (SSC_wire_471, {SSC_wire_471_0, SSC_wire_471_1});
fanout_n #(2, 0, 0) FANOUT_47 (SSC_wire_473, {SSC_wire_473_0, SSC_wire_473_1});
fanout_n #(2, 0, 0) FANOUT_48 (SSC_wire_474, {SSC_wire_474_0, SSC_wire_474_1});
fanout_n #(2, 0, 0) FANOUT_49 (SSC_wire_475, {SSC_wire_475_0, SSC_wire_475_1});
fanout_n #(2, 0, 0) FANOUT_50 (SSC_wire_478, {SSC_wire_478_0, SSC_wire_478_1});
fanout_n #(27, 0, 0) FANOUT_51 (SSC_wire_94, {SSC_wire_94_0, SSC_wire_94_1, SSC_wire_94_2, SSC_wire_94_3, SSC_wire_94_4, SSC_wire_94_5, SSC_wire_94_6, SSC_wire_94_7, SSC_wire_94_8, SSC_wire_94_9, SSC_wire_94_10, SSC_wire_94_11, SSC_wire_94_12, SSC_wire_94_13, SSC_wire_94_14, SSC_wire_94_15, SSC_wire_94_16, SSC_wire_94_17, SSC_wire_94_18, SSC_wire_94_19, SSC_wire_94_20, SSC_wire_94_21, SSC_wire_94_22, SSC_wire_94_23, SSC_wire_94_24, SSC_wire_94_25, SSC_wire_94_26});
fanout_n #(35, 0, 0) FANOUT_52 (SSC_wire_61, {SSC_wire_61_0, SSC_wire_61_1, SSC_wire_61_2, SSC_wire_61_3, SSC_wire_61_4, SSC_wire_61_5, SSC_wire_61_6, SSC_wire_61_7, SSC_wire_61_8, SSC_wire_61_9, SSC_wire_61_10, SSC_wire_61_11, SSC_wire_61_12, SSC_wire_61_13, SSC_wire_61_14, SSC_wire_61_15, SSC_wire_61_16, SSC_wire_61_17, SSC_wire_61_18, SSC_wire_61_19, SSC_wire_61_20, SSC_wire_61_21, SSC_wire_61_22, SSC_wire_61_23, SSC_wire_61_24, SSC_wire_61_25, SSC_wire_61_26, SSC_wire_61_27, SSC_wire_61_28, SSC_wire_61_29, SSC_wire_61_30, SSC_wire_61_31, SSC_wire_61_32, SSC_wire_61_33, SSC_wire_61_34});
fanout_n #(3, 0, 0) FANOUT_53 (SSC_wire_398, {SSC_wire_398_0, SSC_wire_398_1, SSC_wire_398_2});
fanout_n #(28, 0, 0) FANOUT_54 (SSC_wire_20, {SSC_wire_20_0, SSC_wire_20_1, SSC_wire_20_2, SSC_wire_20_3, SSC_wire_20_4, SSC_wire_20_5, SSC_wire_20_6, SSC_wire_20_7, SSC_wire_20_8, SSC_wire_20_9, SSC_wire_20_10, SSC_wire_20_11, SSC_wire_20_12, SSC_wire_20_13, SSC_wire_20_14, SSC_wire_20_15, SSC_wire_20_16, SSC_wire_20_17, SSC_wire_20_18, SSC_wire_20_19, SSC_wire_20_20, SSC_wire_20_21, SSC_wire_20_22, SSC_wire_20_23, SSC_wire_20_24, SSC_wire_20_25, SSC_wire_20_26, SSC_wire_20_27});
fanout_n #(38, 0, 0) FANOUT_55 (SSC_wire_3, {SSC_wire_3_0, SSC_wire_3_1, SSC_wire_3_2, SSC_wire_3_3, SSC_wire_3_4, SSC_wire_3_5, SSC_wire_3_6, SSC_wire_3_7, SSC_wire_3_8, SSC_wire_3_9, SSC_wire_3_10, SSC_wire_3_11, SSC_wire_3_12, SSC_wire_3_13, SSC_wire_3_14, SSC_wire_3_15, SSC_wire_3_16, SSC_wire_3_17, SSC_wire_3_18, SSC_wire_3_19, SSC_wire_3_20, SSC_wire_3_21, SSC_wire_3_22, SSC_wire_3_23, SSC_wire_3_24, SSC_wire_3_25, SSC_wire_3_26, SSC_wire_3_27, SSC_wire_3_28, SSC_wire_3_29, SSC_wire_3_30, SSC_wire_3_31, SSC_wire_3_32, SSC_wire_3_33, SSC_wire_3_34, SSC_wire_3_35, SSC_wire_3_36, SSC_wire_3_37});
fanout_n #(2, 0, 0) FANOUT_56 (SSC_wire_485, {SSC_wire_485_0, SSC_wire_485_1});
fanout_n #(2, 0, 0) FANOUT_57 (SSC_wire_487, {SSC_wire_487_0, SSC_wire_487_1});
fanout_n #(16, 0, 0) FANOUT_58 (SSC_wire_174, {SSC_wire_174_0, SSC_wire_174_1, SSC_wire_174_2, SSC_wire_174_3, SSC_wire_174_4, SSC_wire_174_5, SSC_wire_174_6, SSC_wire_174_7, SSC_wire_174_8, SSC_wire_174_9, SSC_wire_174_10, SSC_wire_174_11, SSC_wire_174_12, SSC_wire_174_13, SSC_wire_174_14, SSC_wire_174_15});
fanout_n #(3, 0, 0) FANOUT_59 (SSC_wire_294, {SSC_wire_294_0, SSC_wire_294_1, SSC_wire_294_2});
fanout_n #(3, 0, 0) FANOUT_60 (SSC_wire_324, {SSC_wire_324_0, SSC_wire_324_1, SSC_wire_324_2});
fanout_n #(3, 0, 0) FANOUT_61 (SSC_wire_322, {SSC_wire_322_0, SSC_wire_322_1, SSC_wire_322_2});
fanout_n #(3, 0, 0) FANOUT_62 (SSC_wire_331, {SSC_wire_331_0, SSC_wire_331_1, SSC_wire_331_2});
fanout_n #(4, 0, 0) FANOUT_63 (SSC_wire_329, {SSC_wire_329_0, SSC_wire_329_1, SSC_wire_329_2, SSC_wire_329_3});
fanout_n #(5, 0, 0) FANOUT_64 (SSC_wire_333, {SSC_wire_333_0, SSC_wire_333_1, SSC_wire_333_2, SSC_wire_333_3, SSC_wire_333_4});
fanout_n #(2, 0, 0) FANOUT_65 (SSC_wire_273, {SSC_wire_273_0, SSC_wire_273_1});
fanout_n #(2, 0, 0) FANOUT_66 (SSC_wire_268, {SSC_wire_268_0, SSC_wire_268_1});
fanout_n #(2, 0, 0) FANOUT_67 (SSC_wire_312, {SSC_wire_312_0, SSC_wire_312_1});
fanout_n #(3, 0, 0) FANOUT_68 (SSC_wire_265, {SSC_wire_265_0, SSC_wire_265_1, SSC_wire_265_2});
fanout_n #(2, 0, 0) FANOUT_69 (SSC_wire_310, {SSC_wire_310_0, SSC_wire_310_1});
fanout_n #(3, 0, 0) FANOUT_70 (SSC_wire_311, {SSC_wire_311_0, SSC_wire_311_1, SSC_wire_311_2});
fanout_n #(3, 0, 0) FANOUT_71 (SSC_wire_318, {SSC_wire_318_0, SSC_wire_318_1, SSC_wire_318_2});
fanout_n #(4, 0, 0) FANOUT_72 (SSC_wire_316, {SSC_wire_316_0, SSC_wire_316_1, SSC_wire_316_2, SSC_wire_316_3});
fanout_n #(2, 0, 0) FANOUT_73 (SSC_wire_307, {SSC_wire_307_0, SSC_wire_307_1});
fanout_n #(8, 0, 0) FANOUT_74 (SSC_wire_399, {SSC_wire_399_0, SSC_wire_399_1, SSC_wire_399_2, SSC_wire_399_3, SSC_wire_399_4, SSC_wire_399_5, SSC_wire_399_6, SSC_wire_399_7});
fanout_n #(3, 0, 0) FANOUT_75 (SSC_wire_504, {SSC_wire_504_0, SSC_wire_504_1, SSC_wire_504_2});


and_n #(2, 0, 0) AND_1 (SSC_wire_1, {SSC_wire_2_0, SSC_wire_3_0});
and_n #(2, 0, 0) AND_2 (SSC_wire_4, {SSC_wire_5_0, SSC_wire_3_1});
and_n #(2, 0, 0) AND_3 (SSC_wire_6, {SSC_wire_7_0, SSC_wire_3_2});
and_n #(2, 0, 0) AND_4 (SSC_wire_8, {SSC_wire_9_0, SSC_wire_3_3});
and_n #(2, 0, 0) AND_5 (SSC_wire_10, {SSC_wire_11_0, SSC_wire_3_4});
and_n #(2, 0, 0) AND_6 (SSC_wire_12, {SSC_wire_13_0, SSC_wire_3_5});
and_n #(2, 0, 0) AND_7 (SSC_wire_14, {SSC_wire_15_0, SSC_wire_3_6});
and_n #(2, 0, 0) AND_8 (SSC_wire_16, {SSC_wire_17_0, SSC_wire_3_7});
and_n #(2, 0, 0) AND_9 (SSC_wire_18, {SSC_wire_19_0, SSC_wire_20_0});
and_n #(2, 0, 0) AND_10 (SSC_wire_21, {SSC_wire_22_0, SSC_wire_20_1});
and_n #(2, 0, 0) AND_11 (SSC_wire_23, {SSC_wire_24_0, SSC_wire_20_2});
and_n #(2, 0, 0) AND_12 (SSC_wire_25, {SSC_wire_26_0, SSC_wire_20_3});
and_n #(2, 0, 0) AND_13 (SSC_wire_27, {SSC_wire_28_0, SSC_wire_20_4});
and_n #(2, 0, 0) AND_14 (SSC_wire_29, {SSC_wire_30_0, SSC_wire_20_5});
and_n #(2, 0, 0) AND_15 (SSC_wire_31, {SSC_wire_32_0, SSC_wire_20_6});
and_n #(2, 0, 0) AND_16 (SSC_wire_33, {SSC_wire_34_0, SSC_wire_20_7});
or_n #(2, 0, 0) OR_1 (SSC_wire_35, {SSC_wire_1, SSC_wire_36});
and_n #(2, 0, 0) AND_17 (SSC_wire_36, {SSC_wire_18, SSC_wire_37});
notg #(0, 0) NOT_1 (SSC_wire_37, SSC_wire_3_8);
or_n #(2, 0, 0) OR_2 (SSC_wire_38, {SSC_wire_4, SSC_wire_39});
and_n #(2, 0, 0) AND_18 (SSC_wire_39, {SSC_wire_21, SSC_wire_40});
notg #(0, 0) NOT_2 (SSC_wire_40, SSC_wire_3_9);
or_n #(2, 0, 0) OR_3 (SSC_wire_41, {SSC_wire_6, SSC_wire_42});
and_n #(2, 0, 0) AND_19 (SSC_wire_42, {SSC_wire_23, SSC_wire_43});
notg #(0, 0) NOT_3 (SSC_wire_43, SSC_wire_3_10);
or_n #(2, 0, 0) OR_4 (SSC_wire_44, {SSC_wire_8, SSC_wire_45});
and_n #(2, 0, 0) AND_20 (SSC_wire_45, {SSC_wire_25, SSC_wire_46});
notg #(0, 0) NOT_4 (SSC_wire_46, SSC_wire_3_11);
or_n #(2, 0, 0) OR_5 (SSC_wire_47, {SSC_wire_10, SSC_wire_48});
and_n #(2, 0, 0) AND_21 (SSC_wire_48, {SSC_wire_27, SSC_wire_49});
notg #(0, 0) NOT_5 (SSC_wire_49, SSC_wire_3_12);
or_n #(2, 0, 0) OR_6 (SSC_wire_50, {SSC_wire_12, SSC_wire_51});
and_n #(2, 0, 0) AND_22 (SSC_wire_51, {SSC_wire_29, SSC_wire_52});
notg #(0, 0) NOT_6 (SSC_wire_52, SSC_wire_3_13);
or_n #(2, 0, 0) OR_7 (SSC_wire_53, {SSC_wire_14, SSC_wire_54});
and_n #(2, 0, 0) AND_23 (SSC_wire_54, {SSC_wire_31, SSC_wire_55});
notg #(0, 0) NOT_7 (SSC_wire_55, SSC_wire_3_14);
or_n #(2, 0, 0) OR_8 (SSC_wire_56, {SSC_wire_16, SSC_wire_57});
and_n #(2, 0, 0) AND_24 (SSC_wire_57, {SSC_wire_33, SSC_wire_58});
notg #(0, 0) NOT_8 (SSC_wire_58, SSC_wire_3_15);
and_n #(2, 0, 0) AND_25 (SSC_wire_59, {SSC_wire_60_0, SSC_wire_61_0});
and_n #(2, 0, 0) AND_26 (SSC_wire_62, {SSC_wire_63_0, SSC_wire_61_1});
and_n #(2, 0, 0) AND_27 (SSC_wire_64, {SSC_wire_65_0, SSC_wire_61_2});
and_n #(2, 0, 0) AND_28 (SSC_wire_66, {SSC_wire_67_0, SSC_wire_61_3});
and_n #(2, 0, 0) AND_29 (SSC_wire_68, {SSC_wire_69_0, SSC_wire_61_4});
and_n #(2, 0, 0) AND_30 (SSC_wire_70, {SSC_wire_71_0, SSC_wire_61_5});
and_n #(2, 0, 0) AND_31 (SSC_wire_72, {SSC_wire_73_0, SSC_wire_61_6});
and_n #(2, 0, 0) AND_32 (SSC_wire_74, {SSC_wire_75_0, SSC_wire_61_7});
and_n #(2, 0, 0) AND_33 (SSC_wire_76, {SSC_wire_77_0, SSC_wire_61_8});
and_n #(2, 0, 0) AND_34 (SSC_wire_78, {SSC_wire_79_0, SSC_wire_61_9});
and_n #(2, 0, 0) AND_35 (SSC_wire_80, {SSC_wire_81_0, SSC_wire_61_10});
and_n #(2, 0, 0) AND_36 (SSC_wire_82, {SSC_wire_83_0, SSC_wire_61_11});
and_n #(2, 0, 0) AND_37 (SSC_wire_84, {SSC_wire_85_0, SSC_wire_61_12});
and_n #(2, 0, 0) AND_38 (SSC_wire_86, {SSC_wire_87_0, SSC_wire_61_13});
and_n #(2, 0, 0) AND_39 (SSC_wire_88, {SSC_wire_89_0, SSC_wire_61_14});
and_n #(2, 0, 0) AND_40 (SSC_wire_90, {SSC_wire_91_0, SSC_wire_61_15});
and_n #(2, 0, 0) AND_41 (SSC_wire_92, {SSC_wire_93, SSC_wire_94_0});
and_n #(2, 0, 0) AND_42 (SSC_wire_95, {SSC_wire_96, SSC_wire_94_1});
and_n #(2, 0, 0) AND_43 (SSC_wire_97, {SSC_wire_98, SSC_wire_94_2});
and_n #(2, 0, 0) AND_44 (SSC_wire_99, {SSC_wire_100, SSC_wire_94_3});
and_n #(2, 0, 0) AND_45 (SSC_wire_101, {SSC_wire_102, SSC_wire_94_4});
and_n #(2, 0, 0) AND_46 (SSC_wire_103, {SSC_wire_104, SSC_wire_94_5});
and_n #(2, 0, 0) AND_47 (SSC_wire_105, {SSC_wire_106, SSC_wire_94_6});
and_n #(2, 0, 0) AND_48 (SSC_wire_107, {SSC_wire_108, SSC_wire_94_7});
and_n #(2, 0, 0) AND_49 (SSC_wire_109, {SSC_wire_110, SSC_wire_94_8});
and_n #(2, 0, 0) AND_50 (SSC_wire_111, {SSC_wire_112, SSC_wire_94_9});
and_n #(2, 0, 0) AND_51 (SSC_wire_113, {SSC_wire_114, SSC_wire_94_10});
and_n #(2, 0, 0) AND_52 (SSC_wire_115, {SSC_wire_116, SSC_wire_94_11});
and_n #(2, 0, 0) AND_53 (SSC_wire_117, {SSC_wire_118, SSC_wire_94_12});
and_n #(2, 0, 0) AND_54 (SSC_wire_119, {SSC_wire_120, SSC_wire_94_13});
and_n #(2, 0, 0) AND_55 (SSC_wire_121, {SSC_wire_122, SSC_wire_94_14});
and_n #(2, 0, 0) AND_56 (SSC_wire_123, {SSC_wire_124, SSC_wire_94_15});
or_n #(2, 0, 0) OR_9 (SSC_wire_125, {SSC_wire_59, SSC_wire_126});
and_n #(2, 0, 0) AND_57 (SSC_wire_126, {SSC_wire_92, SSC_wire_127});
notg #(0, 0) NOT_9 (SSC_wire_127, SSC_wire_61_16);
or_n #(2, 0, 0) OR_10 (SSC_wire_128, {SSC_wire_62, SSC_wire_129});
and_n #(2, 0, 0) AND_58 (SSC_wire_129, {SSC_wire_95, SSC_wire_130});
notg #(0, 0) NOT_10 (SSC_wire_130, SSC_wire_61_17);
or_n #(2, 0, 0) OR_11 (SSC_wire_131, {SSC_wire_64, SSC_wire_132});
and_n #(2, 0, 0) AND_59 (SSC_wire_132, {SSC_wire_97, SSC_wire_133});
notg #(0, 0) NOT_11 (SSC_wire_133, SSC_wire_61_18);
or_n #(2, 0, 0) OR_12 (SSC_wire_134, {SSC_wire_66, SSC_wire_135});
and_n #(2, 0, 0) AND_60 (SSC_wire_135, {SSC_wire_99, SSC_wire_136});
notg #(0, 0) NOT_12 (SSC_wire_136, SSC_wire_61_19);
or_n #(2, 0, 0) OR_13 (SSC_wire_137, {SSC_wire_68, SSC_wire_138});
and_n #(2, 0, 0) AND_61 (SSC_wire_138, {SSC_wire_101, SSC_wire_139});
notg #(0, 0) NOT_13 (SSC_wire_139, SSC_wire_61_20);
or_n #(2, 0, 0) OR_14 (SSC_wire_140, {SSC_wire_70, SSC_wire_141});
and_n #(2, 0, 0) AND_62 (SSC_wire_141, {SSC_wire_103, SSC_wire_142});
notg #(0, 0) NOT_14 (SSC_wire_142, SSC_wire_61_21);
or_n #(2, 0, 0) OR_15 (SSC_wire_143, {SSC_wire_72, SSC_wire_144});
and_n #(2, 0, 0) AND_63 (SSC_wire_144, {SSC_wire_105, SSC_wire_145});
notg #(0, 0) NOT_15 (SSC_wire_145, SSC_wire_61_22);
or_n #(2, 0, 0) OR_16 (SSC_wire_146, {SSC_wire_74, SSC_wire_147});
and_n #(2, 0, 0) AND_64 (SSC_wire_147, {SSC_wire_107, SSC_wire_148});
notg #(0, 0) NOT_16 (SSC_wire_148, SSC_wire_61_23);
or_n #(2, 0, 0) OR_17 (SSC_wire_149, {SSC_wire_76, SSC_wire_150});
and_n #(2, 0, 0) AND_65 (SSC_wire_150, {SSC_wire_109, SSC_wire_151});
notg #(0, 0) NOT_17 (SSC_wire_151, SSC_wire_61_24);
or_n #(2, 0, 0) OR_18 (SSC_wire_152, {SSC_wire_78, SSC_wire_153});
and_n #(2, 0, 0) AND_66 (SSC_wire_153, {SSC_wire_111, SSC_wire_154});
notg #(0, 0) NOT_18 (SSC_wire_154, SSC_wire_61_25);
or_n #(2, 0, 0) OR_19 (SSC_wire_155, {SSC_wire_80, SSC_wire_156});
and_n #(2, 0, 0) AND_67 (SSC_wire_156, {SSC_wire_113, SSC_wire_157});
notg #(0, 0) NOT_19 (SSC_wire_157, SSC_wire_61_26);
or_n #(2, 0, 0) OR_20 (SSC_wire_158, {SSC_wire_82, SSC_wire_159});
and_n #(2, 0, 0) AND_68 (SSC_wire_159, {SSC_wire_115, SSC_wire_160});
notg #(0, 0) NOT_20 (SSC_wire_160, SSC_wire_61_27);
or_n #(2, 0, 0) OR_21 (SSC_wire_161, {SSC_wire_84, SSC_wire_162});
and_n #(2, 0, 0) AND_69 (SSC_wire_162, {SSC_wire_117, SSC_wire_163});
notg #(0, 0) NOT_21 (SSC_wire_163, SSC_wire_61_28);
or_n #(2, 0, 0) OR_22 (SSC_wire_164, {SSC_wire_86, SSC_wire_165});
and_n #(2, 0, 0) AND_70 (SSC_wire_165, {SSC_wire_119, SSC_wire_166});
notg #(0, 0) NOT_22 (SSC_wire_166, SSC_wire_61_29);
or_n #(2, 0, 0) OR_23 (SSC_wire_167, {SSC_wire_88, SSC_wire_168});
and_n #(2, 0, 0) AND_71 (SSC_wire_168, {SSC_wire_121, SSC_wire_169});
notg #(0, 0) NOT_23 (SSC_wire_169, SSC_wire_61_30);
or_n #(2, 0, 0) OR_24 (SSC_wire_170, {SSC_wire_90, SSC_wire_171});
and_n #(2, 0, 0) AND_72 (SSC_wire_171, {SSC_wire_123, SSC_wire_172});
notg #(0, 0) NOT_24 (SSC_wire_172, SSC_wire_61_31);
and_n #(2, 0, 0) AND_73 (SSC_wire_173, {SSC_wire_2_1, SSC_wire_174_0});
and_n #(2, 0, 0) AND_74 (SSC_wire_175, {SSC_wire_5_1, SSC_wire_174_1});
and_n #(2, 0, 0) AND_75 (SSC_wire_176, {SSC_wire_7_1, SSC_wire_174_2});
and_n #(2, 0, 0) AND_76 (SSC_wire_177, {SSC_wire_9_1, SSC_wire_174_3});
and_n #(2, 0, 0) AND_77 (SSC_wire_178, {SSC_wire_11_1, SSC_wire_174_4});
and_n #(2, 0, 0) AND_78 (SSC_wire_179, {SSC_wire_13_1, SSC_wire_174_5});
and_n #(2, 0, 0) AND_79 (SSC_wire_180, {SSC_wire_15_1, SSC_wire_174_6});
and_n #(2, 0, 0) AND_80 (SSC_wire_181, {SSC_wire_17_1, SSC_wire_174_7});
and_n #(2, 0, 0) AND_81 (SSC_wire_182, {SSC_wire_19_1, SSC_wire_20_8});
and_n #(2, 0, 0) AND_82 (SSC_wire_183, {SSC_wire_22_1, SSC_wire_20_9});
and_n #(2, 0, 0) AND_83 (SSC_wire_184, {SSC_wire_24_1, SSC_wire_20_10});
and_n #(2, 0, 0) AND_84 (SSC_wire_185, {SSC_wire_26_1, SSC_wire_20_11});
and_n #(2, 0, 0) AND_85 (SSC_wire_186, {SSC_wire_28_1, SSC_wire_20_12});
and_n #(2, 0, 0) AND_86 (SSC_wire_187, {SSC_wire_30_1, SSC_wire_20_13});
and_n #(2, 0, 0) AND_87 (SSC_wire_188, {SSC_wire_32_1, SSC_wire_20_14});
and_n #(2, 0, 0) AND_88 (SSC_wire_189, {SSC_wire_34_1, SSC_wire_20_15});
and_n #(2, 0, 0) AND_89 (SSC_wire_190, {SSC_wire_191, SSC_wire_94_16});
and_n #(2, 0, 0) AND_90 (SSC_wire_192, {SSC_wire_193, SSC_wire_94_17});
and_n #(2, 0, 0) AND_91 (SSC_wire_194, {SSC_wire_195, SSC_wire_94_18});
and_n #(2, 0, 0) AND_92 (SSC_wire_196, {SSC_wire_197, SSC_wire_94_19});
and_n #(2, 0, 0) AND_93 (SSC_wire_198, {SSC_wire_199, SSC_wire_94_20});
and_n #(2, 0, 0) AND_94 (SSC_wire_200, {SSC_wire_201, SSC_wire_94_21});
and_n #(2, 0, 0) AND_95 (SSC_wire_202, {SSC_wire_203, SSC_wire_94_22});
and_n #(2, 0, 0) AND_96 (SSC_wire_204, {SSC_wire_205, SSC_wire_94_23});
or_n #(2, 0, 0) OR_25 (SSC_wire_206, {SSC_wire_173, SSC_wire_207});
or_n #(2, 0, 0) OR_26 (SSC_wire_208, {SSC_wire_182, SSC_wire_209});
and_n #(2, 0, 0) AND_97 (SSC_wire_209, {SSC_wire_190, SSC_wire_210});
notg #(0, 0) NOT_25 (SSC_wire_210, SSC_wire_20_16);
notg #(0, 0) NOT_26 (SSC_wire_211, SSC_wire_174_8);
and_n #(2, 0, 0) AND_98 (SSC_wire_207, {SSC_wire_211, SSC_wire_208});
or_n #(2, 0, 0) OR_27 (SSC_wire_212, {SSC_wire_175, SSC_wire_213});
or_n #(2, 0, 0) OR_28 (SSC_wire_214, {SSC_wire_183, SSC_wire_215});
and_n #(2, 0, 0) AND_99 (SSC_wire_215, {SSC_wire_192, SSC_wire_216});
notg #(0, 0) NOT_27 (SSC_wire_216, SSC_wire_20_17);
notg #(0, 0) NOT_28 (SSC_wire_217, SSC_wire_174_9);
and_n #(2, 0, 0) AND_100 (SSC_wire_213, {SSC_wire_217, SSC_wire_214});
or_n #(2, 0, 0) OR_29 (SSC_wire_218, {SSC_wire_176, SSC_wire_219});
or_n #(2, 0, 0) OR_30 (SSC_wire_220, {SSC_wire_184, SSC_wire_221});
and_n #(2, 0, 0) AND_101 (SSC_wire_221, {SSC_wire_194, SSC_wire_222});
notg #(0, 0) NOT_29 (SSC_wire_222, SSC_wire_20_18);
notg #(0, 0) NOT_30 (SSC_wire_223, SSC_wire_174_10);
and_n #(2, 0, 0) AND_102 (SSC_wire_219, {SSC_wire_223, SSC_wire_220});
or_n #(2, 0, 0) OR_31 (SSC_wire_224, {SSC_wire_177, SSC_wire_225});
or_n #(2, 0, 0) OR_32 (SSC_wire_226, {SSC_wire_185, SSC_wire_227});
and_n #(2, 0, 0) AND_103 (SSC_wire_227, {SSC_wire_196, SSC_wire_228});
notg #(0, 0) NOT_31 (SSC_wire_228, SSC_wire_20_19);
notg #(0, 0) NOT_32 (SSC_wire_229, SSC_wire_174_11);
and_n #(2, 0, 0) AND_104 (SSC_wire_225, {SSC_wire_229, SSC_wire_226});
or_n #(2, 0, 0) OR_33 (SSC_wire_230, {SSC_wire_178, SSC_wire_231});
or_n #(2, 0, 0) OR_34 (SSC_wire_232, {SSC_wire_186, SSC_wire_233});
and_n #(2, 0, 0) AND_105 (SSC_wire_233, {SSC_wire_198, SSC_wire_234});
notg #(0, 0) NOT_33 (SSC_wire_234, SSC_wire_20_20);
notg #(0, 0) NOT_34 (SSC_wire_235, SSC_wire_174_12);
and_n #(2, 0, 0) AND_106 (SSC_wire_231, {SSC_wire_235, SSC_wire_232});
or_n #(2, 0, 0) OR_35 (SSC_wire_236, {SSC_wire_179, SSC_wire_237});
or_n #(2, 0, 0) OR_36 (SSC_wire_238, {SSC_wire_187, SSC_wire_239});
and_n #(2, 0, 0) AND_107 (SSC_wire_239, {SSC_wire_200, SSC_wire_240});
notg #(0, 0) NOT_35 (SSC_wire_240, SSC_wire_20_21);
notg #(0, 0) NOT_36 (SSC_wire_241, SSC_wire_174_13);
and_n #(2, 0, 0) AND_108 (SSC_wire_237, {SSC_wire_241, SSC_wire_238});
or_n #(2, 0, 0) OR_37 (SSC_wire_242, {SSC_wire_180, SSC_wire_243});
or_n #(2, 0, 0) OR_38 (SSC_wire_244, {SSC_wire_188, SSC_wire_245});
and_n #(2, 0, 0) AND_109 (SSC_wire_245, {SSC_wire_202, SSC_wire_246});
notg #(0, 0) NOT_37 (SSC_wire_246, SSC_wire_20_22);
notg #(0, 0) NOT_38 (SSC_wire_247, SSC_wire_174_14);
and_n #(2, 0, 0) AND_110 (SSC_wire_243, {SSC_wire_247, SSC_wire_244});
or_n #(2, 0, 0) OR_39 (SSC_wire_248, {SSC_wire_181, SSC_wire_249});
or_n #(2, 0, 0) OR_40 (SSC_wire_250, {SSC_wire_189, SSC_wire_251});
and_n #(2, 0, 0) AND_111 (SSC_wire_251, {SSC_wire_204, SSC_wire_252});
notg #(0, 0) NOT_39 (SSC_wire_252, SSC_wire_20_23);
notg #(0, 0) NOT_40 (SSC_wire_253, SSC_wire_174_15);
and_n #(2, 0, 0) AND_112 (SSC_wire_249, {SSC_wire_253, SSC_wire_250});
and_n #(2, 0, 0) AND_113 (SSC_wire_254, {SSC_wire_255, SSC_wire_256});
and_n #(2, 0, 0) AND_114 (SSC_wire_257, {SSC_wire_254, SSC_wire_258});
or_n #(2, 0, 0) OR_41 (SSC_wire_259, {SSC_wire_260, SSC_wire_261});
or_n #(2, 0, 0) OR_42 (SSC_wire_262, {SSC_wire_259, SSC_wire_263});
notg #(0, 0) NOT_41 (SSC_wire_264, SSC_wire_265_0);
or_n #(2, 0, 0) OR_43 (SSC_wire_266, {SSC_wire_264, SSC_wire_81_1});
notg #(0, 0) NOT_42 (SSC_wire_267, SSC_wire_268_0);
and_n #(2, 0, 0) AND_115 (SSC_wire_269, {SSC_wire_267, SSC_wire_77_1});
notg #(0, 0) NOT_43 (SSC_wire_270, SSC_wire_268_1);
or_n #(2, 0, 0) OR_44 (SSC_wire_271, {SSC_wire_270, SSC_wire_77_2});
notg #(0, 0) NOT_44 (SSC_wire_272, SSC_wire_273_0);
and_n #(2, 0, 0) AND_116 (SSC_wire_274, {SSC_wire_272, SSC_wire_75_1});
notg #(0, 0) NOT_45 (SSC_wire_275, SSC_wire_273_1);
or_n #(2, 0, 0) OR_45 (SSC_wire_276, {SSC_wire_275, SSC_wire_75_2});
notg #(0, 0) NOT_46 (SSC_wire_277, SSC_wire_278);
and_n #(3, 0, 0) AND_117 (SSC_wire_279, {SSC_wire_277, SSC_wire_276, SSC_wire_60_1});
notg #(0, 0) NOT_47 (SSC_wire_280, SSC_wire_281);
and_n #(2, 0, 0) AND_118 (SSC_wire_282, {SSC_wire_280, SSC_wire_283});
and_n #(2, 0, 0) AND_119 (SSC_wire_284, {SSC_wire_285, SSC_wire_63_1});
or_n #(2, 0, 0) OR_46 (SSC_wire_263, {SSC_wire_284, SSC_wire_286});
and_n #(2, 0, 0) AND_120 (SSC_wire_286, {SSC_wire_287, SSC_wire_91_1});
and_n #(2, 0, 0) AND_121 (SSC_wire_288, {SSC_wire_289, SSC_wire_81_2});
or_n #(4, 0, 0) OR_47 (SSC_wire_290, {SSC_wire_288, SSC_wire_291, SSC_wire_292, SSC_wire_293});
notg #(0, 0) NOT_48 (SSC_wire_285, SSC_wire_294_0);
and_n #(2, 0, 0) AND_122 (SSC_wire_291, {SSC_wire_295, SSC_wire_83_1});
and_n #(2, 0, 0) AND_123 (SSC_wire_292, {SSC_wire_296, SSC_wire_85_1});
or_n #(2, 0, 0) OR_48 (SSC_wire_297, {SSC_wire_298, SSC_wire_81_3});
and_n #(3, 0, 0) AND_124 (SSC_wire_299, {SSC_wire_297, SSC_wire_300, SSC_wire_79_1});
or_n #(2, 0, 0) OR_49 (SSC_wire_301, {SSC_wire_302, SSC_wire_79_2});
and_n #(2, 0, 0) AND_125 (SSC_wire_303, {SSC_wire_301, SSC_wire_266});
or_n #(2, 0, 0) OR_50 (SSC_wire_304, {SSC_wire_269, SSC_wire_305});
and_n #(2, 0, 0) AND_126 (SSC_wire_305, {SSC_wire_271, SSC_wire_306});
or_n #(2, 0, 0) OR_51 (SSC_wire_306, {SSC_wire_274, SSC_wire_279});
notg #(0, 0) NOT_49 (SSC_wire_287, SSC_wire_307_0);
or_n #(2, 0, 0) OR_52 (SSC_wire_283, {SSC_wire_290, SSC_wire_308});
or_n #(2, 0, 0) OR_53 (SSC_wire_308, {SSC_wire_299, SSC_wire_309});
and_n #(2, 0, 0) AND_127 (SSC_wire_309, {SSC_wire_303, SSC_wire_304});
or_n #(2, 0, 0) OR_54 (SSC_wire_258, {SSC_wire_262, SSC_wire_282});
notg #(0, 0) NOT_50 (SSC_wire_289, SSC_wire_265_1);
notg #(0, 0) NOT_51 (SSC_wire_295, SSC_wire_310_0);
notg #(0, 0) NOT_52 (SSC_wire_296, SSC_wire_311_0);
notg #(0, 0) NOT_53 (SSC_wire_298, SSC_wire_265_2);
notg #(0, 0) NOT_54 (SSC_wire_300, SSC_wire_312_0);
notg #(0, 0) NOT_55 (SSC_wire_302, SSC_wire_312_1);
or_n #(2, 0, 0) OR_55 (SSC_wire_293, {SSC_wire_313, SSC_wire_314});
notg #(0, 0) NOT_56 (SSC_wire_315, SSC_wire_316_0);
and_n #(2, 0, 0) AND_128 (SSC_wire_313, {SSC_wire_315, SSC_wire_89_1});
notg #(0, 0) NOT_57 (SSC_wire_317, SSC_wire_318_0);
and_n #(2, 0, 0) AND_129 (SSC_wire_314, {SSC_wire_317, SSC_wire_87_1});
or_n #(2, 0, 0) OR_56 (SSC_wire_260, {SSC_wire_319, SSC_wire_320});
notg #(0, 0) NOT_58 (SSC_wire_321, SSC_wire_322_0);
and_n #(2, 0, 0) AND_130 (SSC_wire_319, {SSC_wire_321, SSC_wire_67_1});
notg #(0, 0) NOT_59 (SSC_wire_323, SSC_wire_324_0);
and_n #(2, 0, 0) AND_131 (SSC_wire_320, {SSC_wire_323, SSC_wire_65_1});
or_n #(3, 0, 0) OR_57 (SSC_wire_261, {SSC_wire_325, SSC_wire_326, SSC_wire_327});
notg #(0, 0) NOT_60 (SSC_wire_328, SSC_wire_329_0);
and_n #(2, 0, 0) AND_132 (SSC_wire_325, {SSC_wire_328, SSC_wire_71_1});
notg #(0, 0) NOT_61 (SSC_wire_330, SSC_wire_331_0);
and_n #(2, 0, 0) AND_133 (SSC_wire_326, {SSC_wire_330, SSC_wire_69_1});
notg #(0, 0) NOT_62 (SSC_wire_332, SSC_wire_333_0);
and_n #(2, 0, 0) AND_134 (SSC_wire_327, {SSC_wire_332, SSC_wire_73_1});
or_n #(2, 0, 0) OR_58 (SSC_wire_281, {SSC_wire_334, SSC_wire_335});
notg #(0, 0) NOT_63 (SSC_wire_336, SSC_wire_89_2);
and_n #(2, 0, 0) AND_135 (SSC_wire_337, {SSC_wire_336, SSC_wire_316_1});
or_n #(2, 0, 0) OR_59 (SSC_wire_338, {SSC_wire_339, SSC_wire_316_2});
and_n #(3, 0, 0) AND_136 (SSC_wire_340, {SSC_wire_338, SSC_wire_341, SSC_wire_318_1});
or_n #(2, 0, 0) OR_60 (SSC_wire_342, {SSC_wire_343, SSC_wire_316_3});
and_n #(2, 0, 0) AND_137 (SSC_wire_344, {SSC_wire_342, SSC_wire_345});
or_n #(2, 0, 0) OR_61 (SSC_wire_345, {SSC_wire_346, SSC_wire_318_2});
and_n #(2, 0, 0) AND_138 (SSC_wire_347, {SSC_wire_348, SSC_wire_311_1});
or_n #(2, 0, 0) OR_62 (SSC_wire_349, {SSC_wire_347, SSC_wire_350});
or_n #(2, 0, 0) OR_63 (SSC_wire_351, {SSC_wire_352, SSC_wire_311_2});
and_n #(3, 0, 0) AND_139 (SSC_wire_350, {SSC_wire_351, SSC_wire_353, SSC_wire_310_1});
or_n #(2, 0, 0) OR_64 (SSC_wire_334, {SSC_wire_340, SSC_wire_337});
and_n #(2, 0, 0) AND_140 (SSC_wire_335, {SSC_wire_344, SSC_wire_349});
notg #(0, 0) NOT_64 (SSC_wire_339, SSC_wire_89_3);
notg #(0, 0) NOT_65 (SSC_wire_341, SSC_wire_87_2);
notg #(0, 0) NOT_66 (SSC_wire_343, SSC_wire_89_4);
notg #(0, 0) NOT_67 (SSC_wire_346, SSC_wire_87_3);
notg #(0, 0) NOT_68 (SSC_wire_348, SSC_wire_85_2);
notg #(0, 0) NOT_69 (SSC_wire_352, SSC_wire_85_3);
notg #(0, 0) NOT_70 (SSC_wire_353, SSC_wire_83_2);
or_n #(2, 0, 0) OR_65 (SSC_wire_255, {SSC_wire_354, SSC_wire_355});
notg #(0, 0) NOT_71 (SSC_wire_356, SSC_wire_333_1);
and_n #(2, 0, 0) AND_141 (SSC_wire_357, {SSC_wire_356, SSC_wire_73_2});
notg #(0, 0) NOT_72 (SSC_wire_358, SSC_wire_294_1);
and_n #(2, 0, 0) AND_142 (SSC_wire_359, {SSC_wire_358, SSC_wire_63_2});
notg #(0, 0) NOT_73 (SSC_wire_360, SSC_wire_294_2);
or_n #(2, 0, 0) OR_66 (SSC_wire_361, {SSC_wire_360, SSC_wire_63_3});
notg #(0, 0) NOT_74 (SSC_wire_362, SSC_wire_307_1);
or_n #(2, 0, 0) OR_67 (SSC_wire_363, {SSC_wire_362, SSC_wire_91_2});
or_n #(2, 0, 0) OR_68 (SSC_wire_354, {SSC_wire_357, SSC_wire_364});
or_n #(2, 0, 0) OR_69 (SSC_wire_365, {SSC_wire_366, SSC_wire_73_3});
and_n #(2, 0, 0) AND_143 (SSC_wire_364, {SSC_wire_365, SSC_wire_367});
and_n #(2, 0, 0) AND_144 (SSC_wire_368, {SSC_wire_369, SSC_wire_69_2});
or_n #(3, 0, 0) OR_70 (SSC_wire_367, {SSC_wire_368, SSC_wire_370, SSC_wire_371});
and_n #(2, 0, 0) AND_145 (SSC_wire_370, {SSC_wire_372, SSC_wire_67_2});
and_n #(2, 0, 0) AND_146 (SSC_wire_371, {SSC_wire_373, SSC_wire_71_2});
or_n #(2, 0, 0) OR_71 (SSC_wire_374, {SSC_wire_375, SSC_wire_67_3});
and_n #(2, 0, 0) AND_147 (SSC_wire_376, {SSC_wire_374, SSC_wire_377});
or_n #(2, 0, 0) OR_72 (SSC_wire_377, {SSC_wire_378, SSC_wire_73_4});
notg #(0, 0) NOT_75 (SSC_wire_366, SSC_wire_333_2);
and_n #(2, 0, 0) AND_148 (SSC_wire_379, {SSC_wire_380, SSC_wire_65_2});
or_n #(2, 0, 0) OR_73 (SSC_wire_381, {SSC_wire_379, SSC_wire_382});
or_n #(2, 0, 0) OR_74 (SSC_wire_383, {SSC_wire_384, SSC_wire_65_3});
and_n #(2, 0, 0) AND_149 (SSC_wire_382, {SSC_wire_383, SSC_wire_385});
or_n #(2, 0, 0) OR_75 (SSC_wire_385, {SSC_wire_359, SSC_wire_386});
and_n #(2, 0, 0) AND_150 (SSC_wire_386, {SSC_wire_361, SSC_wire_363});
and_n #(2, 0, 0) AND_151 (SSC_wire_355, {SSC_wire_376, SSC_wire_381});
notg #(0, 0) NOT_76 (SSC_wire_369, SSC_wire_331_1);
notg #(0, 0) NOT_77 (SSC_wire_372, SSC_wire_322_1);
notg #(0, 0) NOT_78 (SSC_wire_373, SSC_wire_329_1);
notg #(0, 0) NOT_79 (SSC_wire_375, SSC_wire_322_2);
notg #(0, 0) NOT_80 (SSC_wire_378, SSC_wire_333_3);
notg #(0, 0) NOT_81 (SSC_wire_380, SSC_wire_324_1);
notg #(0, 0) NOT_82 (SSC_wire_384, SSC_wire_324_2);
or_n #(2, 0, 0) OR_76 (SSC_wire_256, {SSC_wire_387, SSC_wire_388});
notg #(0, 0) NOT_83 (SSC_wire_389, SSC_wire_333_4);
and_n #(2, 0, 0) AND_152 (SSC_wire_390, {SSC_wire_389, SSC_wire_73_5});
and_n #(2, 0, 0) AND_153 (SSC_wire_387, {SSC_wire_391, SSC_wire_392});
notg #(0, 0) NOT_84 (SSC_wire_393, SSC_wire_329_2);
and_n #(2, 0, 0) AND_154 (SSC_wire_394, {SSC_wire_393, SSC_wire_71_3});
notg #(0, 0) NOT_85 (SSC_wire_395, SSC_wire_329_3);
or_n #(2, 0, 0) OR_77 (SSC_wire_391, {SSC_wire_395, SSC_wire_71_4});
notg #(0, 0) NOT_86 (SSC_wire_396, SSC_wire_331_2);
or_n #(2, 0, 0) OR_78 (SSC_wire_392, {SSC_wire_396, SSC_wire_69_3});
or_n #(2, 0, 0) OR_79 (SSC_wire_388, {SSC_wire_390, SSC_wire_394});
or_n #(2, 0, 0) OR_80 (SSC_wire_400, {SSC_wire_3_16, SSC_wire_257});
xor_n #(2, 0, 0) XOR_1 (SSC_wire_401, {SSC_wire_402, SSC_wire_34_2});
xor_n #(2, 0, 0) XOR_2 (SSC_wire_403, {SSC_wire_404_0, SSC_wire_32_2});
xor_n #(2, 0, 0) XOR_3 (SSC_wire_405, {SSC_wire_406_0, SSC_wire_30_2});
xor_n #(2, 0, 0) XOR_4 (SSC_wire_407, {SSC_wire_408_0, SSC_wire_28_2});
xor_n #(2, 0, 0) XOR_5 (SSC_wire_409, {SSC_wire_410_0, SSC_wire_26_2});
xor_n #(2, 0, 0) XOR_6 (SSC_wire_411, {SSC_wire_412_0, SSC_wire_24_2});
xor_n #(2, 0, 0) XOR_7 (SSC_wire_413, {SSC_wire_19_2, SSC_wire_22_2});
and_n #(8, 0, 0) AND_155 (SSC_wire_423, {SSC_wire_19_3, SSC_wire_22_3, SSC_wire_24_3, SSC_wire_26_3, SSC_wire_28_3, SSC_wire_30_3, SSC_wire_32_3, SSC_wire_34_3});
and_n #(2, 0, 0) AND_156 (SSC_wire_412, {SSC_wire_19_4, SSC_wire_22_4});
and_n #(2, 0, 0) AND_157 (SSC_wire_410, {SSC_wire_24_4, SSC_wire_412_1});
and_n #(2, 0, 0) AND_158 (SSC_wire_408, {SSC_wire_26_4, SSC_wire_410_1});
and_n #(2, 0, 0) AND_159 (SSC_wire_406, {SSC_wire_28_4, SSC_wire_408_1});
and_n #(2, 0, 0) AND_160 (SSC_wire_404, {SSC_wire_30_4, SSC_wire_406_1});
and_n #(2, 0, 0) AND_161 (SSC_wire_402, {SSC_wire_32_4, SSC_wire_404_1});
or_n #(2, 0, 0) OR_81 (SSC_wire_415, {SSC_wire_424, SSC_wire_425});
and_n #(2, 0, 0) AND_162 (SSC_wire_424, {SSC_wire_3_17, SSC_wire_426});
nor_n #(2, 0, 0) NOR_1 (SSC_wire_425, {SSC_wire_3_18, SSC_wire_19_5});
or_n #(2, 0, 0) OR_82 (SSC_wire_416, {SSC_wire_427, SSC_wire_428});
and_n #(2, 0, 0) AND_163 (SSC_wire_427, {SSC_wire_3_19, SSC_wire_429});
notg #(0, 0) NOT_87 (SSC_wire_430, SSC_wire_3_20);
and_n #(2, 0, 0) AND_164 (SSC_wire_428, {SSC_wire_430, SSC_wire_413});
or_n #(2, 0, 0) OR_83 (SSC_wire_417, {SSC_wire_431, SSC_wire_432});
and_n #(2, 0, 0) AND_165 (SSC_wire_431, {SSC_wire_3_21, SSC_wire_433});
notg #(0, 0) NOT_88 (SSC_wire_434, SSC_wire_3_22);
and_n #(2, 0, 0) AND_166 (SSC_wire_432, {SSC_wire_434, SSC_wire_411});
or_n #(2, 0, 0) OR_84 (SSC_wire_418, {SSC_wire_435, SSC_wire_436});
and_n #(2, 0, 0) AND_167 (SSC_wire_435, {SSC_wire_3_23, SSC_wire_437});
notg #(0, 0) NOT_89 (SSC_wire_438, SSC_wire_3_24);
and_n #(2, 0, 0) AND_168 (SSC_wire_436, {SSC_wire_438, SSC_wire_409});
or_n #(2, 0, 0) OR_85 (SSC_wire_419, {SSC_wire_439, SSC_wire_440});
and_n #(2, 0, 0) AND_169 (SSC_wire_439, {SSC_wire_3_25, SSC_wire_441});
notg #(0, 0) NOT_90 (SSC_wire_442, SSC_wire_3_26);
and_n #(2, 0, 0) AND_170 (SSC_wire_440, {SSC_wire_442, SSC_wire_407});
or_n #(2, 0, 0) OR_86 (SSC_wire_420, {SSC_wire_443, SSC_wire_444});
and_n #(2, 0, 0) AND_171 (SSC_wire_443, {SSC_wire_3_27, SSC_wire_445});
notg #(0, 0) NOT_91 (SSC_wire_446, SSC_wire_3_28);
and_n #(2, 0, 0) AND_172 (SSC_wire_444, {SSC_wire_446, SSC_wire_405});
or_n #(2, 0, 0) OR_87 (SSC_wire_421, {SSC_wire_447, SSC_wire_448});
and_n #(2, 0, 0) AND_173 (SSC_wire_447, {SSC_wire_3_29, SSC_wire_449});
notg #(0, 0) NOT_92 (SSC_wire_450, SSC_wire_3_30);
and_n #(2, 0, 0) AND_174 (SSC_wire_448, {SSC_wire_450, SSC_wire_403});
or_n #(2, 0, 0) OR_88 (SSC_wire_422, {SSC_wire_451, SSC_wire_452});
and_n #(2, 0, 0) AND_175 (SSC_wire_451, {SSC_wire_3_31, SSC_wire_453});
notg #(0, 0) NOT_93 (SSC_wire_454, SSC_wire_3_32);
and_n #(2, 0, 0) AND_176 (SSC_wire_452, {SSC_wire_454, SSC_wire_401});
or_n #(2, 0, 0) OR_89 (SSC_wire_414, {SSC_wire_455, SSC_wire_3_33});
xor_n #(2, 0, 0) XOR_8 (SSC_wire_456, {SSC_wire_457, SSC_wire_17_2});
xor_n #(2, 0, 0) XOR_9 (SSC_wire_458, {SSC_wire_459_0, SSC_wire_15_2});
xor_n #(2, 0, 0) XOR_10 (SSC_wire_460, {SSC_wire_461_0, SSC_wire_13_2});
xor_n #(2, 0, 0) XOR_11 (SSC_wire_462, {SSC_wire_463_0, SSC_wire_11_2});
xor_n #(2, 0, 0) XOR_12 (SSC_wire_464, {SSC_wire_465_0, SSC_wire_9_2});
xor_n #(2, 0, 0) XOR_13 (SSC_wire_466, {SSC_wire_467_0, SSC_wire_7_2});
xor_n #(2, 0, 0) XOR_14 (SSC_wire_468, {SSC_wire_2_2, SSC_wire_5_2});
and_n #(8, 0, 0) AND_177 (SSC_wire_470, {SSC_wire_2_3, SSC_wire_5_3, SSC_wire_7_3, SSC_wire_9_3, SSC_wire_11_3, SSC_wire_13_3, SSC_wire_15_3, SSC_wire_17_3});
notg #(0, 0) NOT_94 (SSC_wire_469, SSC_wire_2_4);
and_n #(2, 0, 0) AND_178 (SSC_wire_467, {SSC_wire_2_5, SSC_wire_5_4});
and_n #(2, 0, 0) AND_179 (SSC_wire_465, {SSC_wire_7_4, SSC_wire_467_1});
and_n #(2, 0, 0) AND_180 (SSC_wire_463, {SSC_wire_9_4, SSC_wire_465_1});
and_n #(2, 0, 0) AND_181 (SSC_wire_461, {SSC_wire_11_4, SSC_wire_463_1});
and_n #(2, 0, 0) AND_182 (SSC_wire_459, {SSC_wire_13_4, SSC_wire_461_1});
and_n #(2, 0, 0) AND_183 (SSC_wire_457, {SSC_wire_15_4, SSC_wire_459_1});
xor_n #(2, 0, 0) XOR_15 (SSC_wire_429, {SSC_wire_2_6, SSC_wire_5_5});
xor_n #(2, 0, 0) XOR_16 (SSC_wire_433, {SSC_wire_471_0, SSC_wire_7_5});
xor_n #(2, 0, 0) XOR_17 (SSC_wire_437, {SSC_wire_472_0, SSC_wire_9_5});
xor_n #(2, 0, 0) XOR_18 (SSC_wire_441, {SSC_wire_473_0, SSC_wire_11_5});
xor_n #(2, 0, 0) XOR_19 (SSC_wire_445, {SSC_wire_474_0, SSC_wire_13_5});
xor_n #(2, 0, 0) XOR_20 (SSC_wire_449, {SSC_wire_475_0, SSC_wire_15_5});
xor_n #(2, 0, 0) XOR_21 (SSC_wire_453, {SSC_wire_476, SSC_wire_17_4});
and_n #(2, 0, 0) AND_184 (SSC_wire_472, {SSC_wire_471_1, SSC_wire_7_6});
and_n #(2, 0, 0) AND_185 (SSC_wire_471, {SSC_wire_2_7, SSC_wire_5_6});
and_n #(2, 0, 0) AND_186 (SSC_wire_473, {SSC_wire_472_1, SSC_wire_9_6});
and_n #(2, 0, 0) AND_187 (SSC_wire_474, {SSC_wire_473_1, SSC_wire_11_6});
and_n #(2, 0, 0) AND_188 (SSC_wire_475, {SSC_wire_474_1, SSC_wire_13_6});
and_n #(2, 0, 0) AND_189 (SSC_wire_476, {SSC_wire_475_1, SSC_wire_15_6});
notg #(0, 0) NOT_95 (SSC_wire_426, SSC_wire_2_8);
and_n #(2, 0, 0) AND_190 (SSC_wire_488, {SSC_wire_470_0, SSC_wire_94_24});
notg #(0, 0) NOT_96 (SSC_wire_489, SSC_wire_470_1);
notg #(0, 0) NOT_97 (SSC_wire_490, SSC_wire_423_0);
and_n #(2, 0, 0) AND_191 (SSC_wire_491, {SSC_wire_423_1, SSC_wire_20_24});
or_n #(2, 0, 0) OR_90 (SSC_wire_455, {SSC_wire_20_25, SSC_wire_3_34});
or_n #(2, 0, 0) OR_91 (SSC_wire_492, {SSC_wire_478_0, SSC_wire_399_0});
and_n #(2, 0, 0) AND_192 (SSC_wire_477, {SSC_wire_488, SSC_wire_493});
notg #(0, 0) NOT_98 (SSC_wire_493, SSC_wire_399_1);
or_n #(2, 0, 0) OR_92 (SSC_wire_494, {SSC_wire_94_25, SSC_wire_61_32});
and_n #(2, 0, 0) AND_193 (SSC_wire_495, {SSC_wire_94_26, SSC_wire_489});
notg #(0, 0) NOT_99 (SSC_wire_496, SSC_wire_399_2);
and_n #(2, 0, 0) AND_194 (SSC_wire_479, {SSC_wire_496, SSC_wire_61_33});
or_n #(3, 0, 0) OR_93 (SSC_wire_174, {SSC_wire_61_34, SSC_wire_398_0, SSC_wire_3_35});
notg #(0, 0) NOT_100 (SSC_wire_497, SSC_wire_399_3);
and_n #(2, 0, 0) AND_195 (SSC_wire_480, {SSC_wire_497, SSC_wire_398_1});
or_n #(3, 0, 0) OR_94 (SSC_wire_498, {SSC_wire_398_2, SSC_wire_20_26, SSC_wire_3_36});
and_n #(2, 0, 0) AND_196 (SSC_wire_481, {SSC_wire_491, SSC_wire_499});
notg #(0, 0) NOT_101 (SSC_wire_499, SSC_wire_399_4);
and_n #(2, 0, 0) AND_197 (SSC_wire_500, {SSC_wire_20_27, SSC_wire_490});
notg #(0, 0) NOT_102 (SSC_wire_501, SSC_wire_399_5);
and_n #(2, 0, 0) AND_198 (SSC_wire_482, {SSC_wire_501, SSC_wire_502});
or_n #(2, 0, 0) OR_95 (SSC_wire_502, {SSC_wire_500, SSC_wire_3_37});
notg #(0, 0) NOT_103 (SSC_wire_503, SSC_wire_504_0);
and_n #(2, 0, 0) AND_199 (SSC_wire_505, {SSC_wire_503, SSC_wire_485_0});
notg #(0, 0) NOT_104 (SSC_wire_506, SSC_wire_399_6);
and_n #(2, 0, 0) AND_200 (SSC_wire_483, {SSC_wire_506, SSC_wire_507});
or_n #(2, 0, 0) OR_96 (SSC_wire_507, {SSC_wire_505, SSC_wire_495});
or_n #(2, 0, 0) OR_97 (SSC_wire_508, {SSC_wire_485_1, SSC_wire_487_0});
and_n #(3, 0, 0) AND_201 (SSC_wire_484, {SSC_wire_508, SSC_wire_509, SSC_wire_504_1});
notg #(0, 0) NOT_105 (SSC_wire_509, SSC_wire_399_7);
and_n #(2, 0, 0) AND_202 (SSC_wire_510, {SSC_wire_487_1, SSC_wire_511});
or_n #(2, 0, 0) OR_98 (SSC_wire_486, {SSC_wire_492, SSC_wire_510});
notg #(0, 0) NOT_106 (SSC_wire_511, SSC_wire_504_2);
bufg #(0, 0) BUF_1 (addr_7, SSC_wire_206);
bufg #(0, 0) BUF_2 (addr_6, SSC_wire_212);
bufg #(0, 0) BUF_3 (addr_5, SSC_wire_218);
bufg #(0, 0) BUF_4 (addr_4, SSC_wire_224);
bufg #(0, 0) BUF_5 (addr_3, SSC_wire_230);
bufg #(0, 0) BUF_6 (addr_2, SSC_wire_236);
bufg #(0, 0) BUF_7 (addr_1, SSC_wire_242);
bufg #(0, 0) BUF_8 (addr_0, SSC_wire_248);
bufg #(0, 0) BUF_9 (SSC_wire_397, clk_net_0);
bufg #(0, 0) BUF_10 (done_net_0, SSC_wire_478_1);
bufg #(0, 0) BUF_11 (read_reg_net_0, SSC_wire_498);
bufg #(0, 0) BUF_12 (SSC_wire_278, readdata_15);
bufg #(0, 0) BUF_13 (SSC_wire_294, readdata_5);
bufg #(0, 0) BUF_14 (SSC_wire_324, readdata_4);
bufg #(0, 0) BUF_15 (SSC_wire_322, readdata_3);
bufg #(0, 0) BUF_16 (SSC_wire_331, readdata_2);
bufg #(0, 0) BUF_17 (SSC_wire_329, readdata_1);
bufg #(0, 0) BUF_18 (SSC_wire_333, readdata_0);
bufg #(0, 0) BUF_19 (SSC_wire_273, readdata_14);
bufg #(0, 0) BUF_20 (SSC_wire_268, readdata_13);
bufg #(0, 0) BUF_21 (SSC_wire_312, readdata_12);
bufg #(0, 0) BUF_22 (SSC_wire_265, readdata_11);
bufg #(0, 0) BUF_23 (SSC_wire_310, readdata_10);
bufg #(0, 0) BUF_24 (SSC_wire_311, readdata_9);
bufg #(0, 0) BUF_25 (SSC_wire_318, readdata_8);
bufg #(0, 0) BUF_26 (SSC_wire_316, readdata_7);
bufg #(0, 0) BUF_27 (SSC_wire_307, readdata_6);
bufg #(0, 0) BUF_28 (SSC_wire_399, rst_net_0);
bufg #(0, 0) BUF_29 (SSC_wire_504, start_net_0);
bufg #(0, 0) BUF_30 (write_reg_net_0, SSC_wire_494);
bufg #(0, 0) BUF_31 (writedata_15, SSC_wire_125);
bufg #(0, 0) BUF_32 (writedata_5, SSC_wire_128);
bufg #(0, 0) BUF_33 (writedata_4, SSC_wire_131);
bufg #(0, 0) BUF_34 (writedata_3, SSC_wire_134);
bufg #(0, 0) BUF_35 (writedata_2, SSC_wire_137);
bufg #(0, 0) BUF_36 (writedata_1, SSC_wire_140);
bufg #(0, 0) BUF_37 (writedata_0, SSC_wire_143);
bufg #(0, 0) BUF_38 (writedata_14, SSC_wire_146);
bufg #(0, 0) BUF_39 (writedata_13, SSC_wire_149);
bufg #(0, 0) BUF_40 (writedata_12, SSC_wire_152);
bufg #(0, 0) BUF_41 (writedata_11, SSC_wire_155);
bufg #(0, 0) BUF_42 (writedata_10, SSC_wire_158);
bufg #(0, 0) BUF_43 (writedata_9, SSC_wire_161);
bufg #(0, 0) BUF_44 (writedata_8, SSC_wire_164);
bufg #(0, 0) BUF_45 (writedata_7, SSC_wire_167);
bufg #(0, 0) BUF_46 (writedata_6, SSC_wire_170);
dff DFF_1  (SSC_wire_106, SSC_wire_333, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_398, NbarT, Si, 1'b0);
dff DFF_2  (SSC_wire_104, SSC_wire_329, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_398, NbarT, SSC_wire_106, 1'b0);
dff DFF_3  (SSC_wire_102, SSC_wire_331, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_398, NbarT, SSC_wire_104, 1'b0);
dff DFF_4  (SSC_wire_100, SSC_wire_322, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_398, NbarT, SSC_wire_102, 1'b0);
dff DFF_5  (SSC_wire_98, SSC_wire_324, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_398, NbarT, SSC_wire_100, 1'b0);
dff DFF_6  (SSC_wire_96, SSC_wire_294, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_398, NbarT, SSC_wire_98, 1'b0);
dff DFF_7  (SSC_wire_124, SSC_wire_307, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_398, NbarT, SSC_wire_96, 1'b0);
dff DFF_8  (SSC_wire_122, SSC_wire_316, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_398, NbarT, SSC_wire_124, 1'b0);
dff DFF_9  (SSC_wire_120, SSC_wire_318, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_398, NbarT, SSC_wire_122, 1'b0);
dff DFF_10  (SSC_wire_118, SSC_wire_311, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_398, NbarT, SSC_wire_120, 1'b0);
dff DFF_11  (SSC_wire_116, SSC_wire_310, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_398, NbarT, SSC_wire_118, 1'b0);
dff DFF_12  (SSC_wire_114, SSC_wire_265, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_398, NbarT, SSC_wire_116, 1'b0);
dff DFF_13  (SSC_wire_112, SSC_wire_312, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_398, NbarT, SSC_wire_114, 1'b0);
dff DFF_14  (SSC_wire_110, SSC_wire_268, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_398, NbarT, SSC_wire_112, 1'b0);
dff DFF_15  (SSC_wire_108, SSC_wire_273, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_398, NbarT, SSC_wire_110, 1'b0);
dff DFF_16  (SSC_wire_93, SSC_wire_278, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_398, NbarT, SSC_wire_108, 1'b0);
dff DFF_17  (SSC_wire_73, SSC_wire_333, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_93, 1'b0);
dff DFF_18  (SSC_wire_71, SSC_wire_329, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_73, 1'b0);
dff DFF_19  (SSC_wire_69, SSC_wire_331, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_71, 1'b0);
dff DFF_20  (SSC_wire_67, SSC_wire_322, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_69, 1'b0);
dff DFF_21  (SSC_wire_65, SSC_wire_324, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_67, 1'b0);
dff DFF_22  (SSC_wire_63, SSC_wire_294, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_65, 1'b0);
dff DFF_23  (SSC_wire_91, SSC_wire_307, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_63, 1'b0);
dff DFF_24  (SSC_wire_89, SSC_wire_316, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_91, 1'b0);
dff DFF_25  (SSC_wire_87, SSC_wire_318, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_89, 1'b0);
dff DFF_26  (SSC_wire_85, SSC_wire_311, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_87, 1'b0);
dff DFF_27  (SSC_wire_83, SSC_wire_310, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_85, 1'b0);
dff DFF_28  (SSC_wire_81, SSC_wire_265, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_83, 1'b0);
dff DFF_29  (SSC_wire_79, SSC_wire_312, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_81, 1'b0);
dff DFF_30  (SSC_wire_77, SSC_wire_268, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_79, 1'b0);
dff DFF_31  (SSC_wire_75, SSC_wire_273, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_77, 1'b0);
dff DFF_32  (SSC_wire_60, SSC_wire_278, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_75, 1'b0);
dff DFF_33  (SSC_wire_205, SSC_wire_56, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_60, 1'b0);
dff DFF_34  (SSC_wire_203, SSC_wire_53, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_205, 1'b0);
dff DFF_35  (SSC_wire_201, SSC_wire_50, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_203, 1'b0);
dff DFF_36  (SSC_wire_199, SSC_wire_47, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_201, 1'b0);
dff DFF_37  (SSC_wire_197, SSC_wire_44, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_199, 1'b0);
dff DFF_38  (SSC_wire_195, SSC_wire_41, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_197, 1'b0);
dff DFF_39  (SSC_wire_193, SSC_wire_38, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_195, 1'b0);
dff DFF_40  (SSC_wire_191, SSC_wire_35, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_400, NbarT, SSC_wire_193, 1'b0);
dff DFF_41  (SSC_wire_19, SSC_wire_415, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_414, NbarT, SSC_wire_191, 1'b0);
dff DFF_42  (SSC_wire_22, SSC_wire_416, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_414, NbarT, SSC_wire_19, 1'b0);
dff DFF_43  (SSC_wire_24, SSC_wire_417, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_414, NbarT, SSC_wire_22, 1'b0);
dff DFF_44  (SSC_wire_26, SSC_wire_418, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_414, NbarT, SSC_wire_24, 1'b0);
dff DFF_45  (SSC_wire_28, SSC_wire_419, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_414, NbarT, SSC_wire_26, 1'b0);
dff DFF_46  (SSC_wire_30, SSC_wire_420, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_414, NbarT, SSC_wire_28, 1'b0);
dff DFF_47  (SSC_wire_32, SSC_wire_421, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_414, NbarT, SSC_wire_30, 1'b0);
dff DFF_48  (SSC_wire_34, SSC_wire_422, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_414, NbarT, SSC_wire_32, 1'b0);
dff DFF_49  (SSC_wire_2, SSC_wire_469, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_61, NbarT, SSC_wire_34, 1'b0);
dff DFF_50  (SSC_wire_5, SSC_wire_468, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_61, NbarT, SSC_wire_2, 1'b0);
dff DFF_51  (SSC_wire_7, SSC_wire_466, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_61, NbarT, SSC_wire_5, 1'b0);
dff DFF_52  (SSC_wire_9, SSC_wire_464, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_61, NbarT, SSC_wire_7, 1'b0);
dff DFF_53  (SSC_wire_11, SSC_wire_462, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_61, NbarT, SSC_wire_9, 1'b0);
dff DFF_54  (SSC_wire_13, SSC_wire_460, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_61, NbarT, SSC_wire_11, 1'b0);
dff DFF_55  (SSC_wire_15, SSC_wire_458, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_61, NbarT, SSC_wire_13, 1'b0);
dff DFF_56  (SSC_wire_17, SSC_wire_456, SSC_wire_397, SSC_wire_399, 1'b0, SSC_wire_61, NbarT, SSC_wire_15, 1'b0);
dff DFF_57  (SSC_wire_478, SSC_wire_477, SSC_wire_397, 1'b0, 1'b0, 1'b1, NbarT, SSC_wire_17, 1'b0);
dff DFF_58  (SSC_wire_94, SSC_wire_479, SSC_wire_397, 1'b0, 1'b0, 1'b1, NbarT, SSC_wire_478, 1'b0);
dff DFF_59  (SSC_wire_61, SSC_wire_480, SSC_wire_397, 1'b0, 1'b0, 1'b1, NbarT, SSC_wire_94, 1'b0);
dff DFF_60  (SSC_wire_398, SSC_wire_481, SSC_wire_397, 1'b0, 1'b0, 1'b1, NbarT, SSC_wire_61, 1'b0);
dff DFF_61  (SSC_wire_20, SSC_wire_482, SSC_wire_397, 1'b0, 1'b0, 1'b1, NbarT, SSC_wire_398, 1'b0);
dff DFF_62  (SSC_wire_3, SSC_wire_483, SSC_wire_397, 1'b0, 1'b0, 1'b1, NbarT, SSC_wire_20, 1'b0);
dff DFF_63  (SSC_wire_485, SSC_wire_484, SSC_wire_397, 1'b0, 1'b0, 1'b1, NbarT, SSC_wire_3, 1'b0);
dff DFF_64  (SSC_wire_487, SSC_wire_486, SSC_wire_397, 1'b0, 1'b0, 1'b1, NbarT, SSC_wire_485, 1'b0);

assign So = SSC_wire_487;

endmodule
